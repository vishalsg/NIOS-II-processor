
module nios_2_DW01_add_8 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267;

  CND3X2 U2 ( .A(n102), .B(n103), .C(n104), .Z(n101) );
  COND3X1 U3 ( .A(n98), .B(n99), .C(n100), .D(n101), .Z(n1) );
  COR2X1 U4 ( .A(B[8]), .B(A[8]), .Z(n25) );
  CND2XL U5 ( .A(n21), .B(n25), .Z(n252) );
  CIVXL U6 ( .A(n25), .Z(n18) );
  CENXL U7 ( .A(n94), .B(n95), .Z(SUM[26]) );
  CIVXL U8 ( .A(n218), .Z(n224) );
  COND1XL U9 ( .A(n112), .B(n113), .C(n114), .Z(n108) );
  CAN2XL U10 ( .A(n265), .B(n142), .Z(SUM[0]) );
  CAN2X1 U11 ( .A(n42), .B(n43), .Z(n3) );
  CAN2X1 U12 ( .A(n180), .B(n181), .Z(n4) );
  CAN2X1 U13 ( .A(n107), .B(n108), .Z(n5) );
  CND2X1 U14 ( .A(B[14]), .B(A[14]), .Z(n198) );
  COR2X1 U15 ( .A(B[14]), .B(A[14]), .Z(n211) );
  COND1X1 U16 ( .A(n37), .B(n3), .C(n38), .Z(n33) );
  CND2XL U17 ( .A(n173), .B(n175), .Z(n248) );
  CND2XL U18 ( .A(n39), .B(n44), .Z(n258) );
  CND2XL U19 ( .A(n44), .B(n42), .Z(n45) );
  CND2XL U20 ( .A(n44), .B(n27), .Z(n43) );
  CND2XL U21 ( .A(n42), .B(n38), .Z(n185) );
  CIVX1 U22 ( .A(n246), .Z(n171) );
  CND2XL U23 ( .A(n175), .B(n234), .Z(n244) );
  CND2XL U24 ( .A(n234), .B(n250), .Z(n249) );
  CND2X2 U25 ( .A(n162), .B(n163), .Z(n104) );
  CNR2X2 U26 ( .A(n186), .B(n187), .Z(n162) );
  COR2X1 U27 ( .A(B[26]), .B(A[26]), .Z(n93) );
  CENXL U28 ( .A(n97), .B(n1), .Z(SUM[25]) );
  CND2X1 U29 ( .A(B[15]), .B(A[15]), .Z(n197) );
  COR2X1 U30 ( .A(B[15]), .B(A[15]), .Z(n193) );
  CND2X1 U31 ( .A(B[5]), .B(A[5]), .Z(n38) );
  COR2X1 U32 ( .A(B[5]), .B(A[5]), .Z(n39) );
  COR2X1 U33 ( .A(B[27]), .B(A[27]), .Z(n86) );
  COR2X1 U34 ( .A(B[17]), .B(A[17]), .Z(n155) );
  COR2X1 U35 ( .A(B[20]), .B(A[20]), .Z(n130) );
  CIVXL U36 ( .A(B[0]), .Z(n266) );
  CND2X2 U37 ( .A(B[0]), .B(A[0]), .Z(n142) );
  CND2X1 U38 ( .A(B[7]), .B(A[7]), .Z(n32) );
  COR2X1 U39 ( .A(B[7]), .B(A[7]), .Z(n31) );
  CND2X1 U40 ( .A(B[10]), .B(A[10]), .Z(n174) );
  COR2X1 U41 ( .A(B[10]), .B(A[10]), .Z(n234) );
  CND2X1 U42 ( .A(B[3]), .B(A[3]), .Z(n48) );
  COR2X1 U43 ( .A(B[3]), .B(A[3]), .Z(n49) );
  CND2X1 U44 ( .A(B[21]), .B(A[21]), .Z(n128) );
  COR2X1 U45 ( .A(B[21]), .B(A[21]), .Z(n129) );
  CND2X1 U46 ( .A(B[2]), .B(A[2]), .Z(n73) );
  COR2X1 U47 ( .A(B[2]), .B(A[2]), .Z(n51) );
  CND2X1 U48 ( .A(B[6]), .B(A[6]), .Z(n40) );
  COR2X1 U49 ( .A(B[6]), .B(A[6]), .Z(n34) );
  CND2X1 U50 ( .A(B[12]), .B(A[12]), .Z(n221) );
  COR2X1 U51 ( .A(B[12]), .B(A[12]), .Z(n233) );
  COR2X1 U52 ( .A(B[11]), .B(A[11]), .Z(n175) );
  CND2X1 U53 ( .A(B[9]), .B(A[9]), .Z(n22) );
  COR2X1 U54 ( .A(B[9]), .B(A[9]), .Z(n21) );
  CIVXL U55 ( .A(n149), .Z(n147) );
  CNR2X1 U56 ( .A(n176), .B(n207), .Z(n205) );
  CND2XL U57 ( .A(n175), .B(n233), .Z(n232) );
  CENXL U58 ( .A(n74), .B(n75), .Z(SUM[29]) );
  CNR2IX1 U59 ( .B(n198), .A(n216), .Z(n214) );
  COND1XL U60 ( .A(n146), .B(n147), .C(n148), .Z(n138) );
  CNR2IXL U61 ( .B(n193), .A(n194), .Z(n188) );
  CNR2XL U62 ( .A(n253), .B(n28), .Z(n19) );
  CNR2XL U63 ( .A(n241), .B(n178), .Z(n253) );
  CNR2XL U64 ( .A(n178), .B(n179), .Z(n191) );
  CND2XL U65 ( .A(n203), .B(n204), .Z(n202) );
  CNR2IXL U66 ( .B(n84), .A(n82), .Z(n88) );
  COND1X1 U67 ( .A(n89), .B(n90), .C(n91), .Z(n85) );
  COND4CXL U68 ( .A(n171), .B(n172), .C(n245), .D(n175), .Z(n231) );
  CND2XL U69 ( .A(n173), .B(n174), .Z(n245) );
  COND4CXL U70 ( .A(n26), .B(n27), .C(n228), .D(n229), .Z(n218) );
  CND2XL U71 ( .A(n207), .B(n192), .Z(n261) );
  CND2XL U72 ( .A(n51), .B(n73), .Z(n68) );
  CEOXL U73 ( .A(n151), .B(n152), .Z(SUM[18]) );
  CEOXL U74 ( .A(n144), .B(n145), .Z(SUM[19]) );
  CEOXL U75 ( .A(n124), .B(n125), .Z(SUM[22]) );
  CEOXL U76 ( .A(n109), .B(n110), .Z(SUM[24]) );
  CEOXL U77 ( .A(n117), .B(n118), .Z(SUM[23]) );
  CEOXL U78 ( .A(n134), .B(n135), .Z(SUM[20]) );
  CND2XL U79 ( .A(n130), .B(n127), .Z(n135) );
  CNR2IXL U80 ( .B(n221), .A(n224), .Z(n226) );
  CEOXL U81 ( .A(n29), .B(n30), .Z(SUM[7]) );
  CND2XL U82 ( .A(n31), .B(n32), .Z(n30) );
  CNR2IXL U83 ( .B(n32), .A(n14), .Z(n254) );
  CND2XL U84 ( .A(n234), .B(n174), .Z(n251) );
  CND2XL U85 ( .A(n92), .B(n90), .Z(n97) );
  CNR2XL U86 ( .A(n48), .B(n176), .Z(n203) );
  CNR2IXL U87 ( .B(n175), .A(n176), .Z(n167) );
  CND3XL U88 ( .A(n49), .B(n262), .C(n263), .Z(n207) );
  CND2XL U89 ( .A(n21), .B(n22), .Z(n16) );
  CND2XL U90 ( .A(n48), .B(n49), .Z(n47) );
  CND2XL U91 ( .A(n155), .B(n153), .Z(n158) );
  CEOXL U92 ( .A(n157), .B(n158), .Z(SUM[17]) );
  CENXL U93 ( .A(n247), .B(n248), .Z(SUM[11]) );
  CANR4CXL U94 ( .A(n177), .B(n224), .C(n220), .D(n225), .Z(n222) );
  CEOXL U95 ( .A(n222), .B(n223), .Z(SUM[14]) );
  CND2XL U96 ( .A(n211), .B(n198), .Z(n223) );
  CND2XL U97 ( .A(n173), .B(n174), .Z(n169) );
  CNR2XL U98 ( .A(n195), .B(n196), .Z(n194) );
  COND1X1 U99 ( .A(n119), .B(n120), .C(n121), .Z(n115) );
  CIVXL U100 ( .A(n122), .Z(n120) );
  CIVXL U101 ( .A(n115), .Z(n113) );
  CENXL U102 ( .A(n36), .B(n33), .Z(SUM[6]) );
  CENX1 U103 ( .A(n53), .B(n54), .Z(SUM[31]) );
  CND2XL U104 ( .A(B[8]), .B(A[8]), .Z(n20) );
  CND2XL U105 ( .A(B[4]), .B(A[4]), .Z(n42) );
  COR2XL U106 ( .A(B[13]), .B(A[13]), .Z(n220) );
  CND2XL U107 ( .A(B[1]), .B(A[1]), .Z(n71) );
  COR2XL U108 ( .A(B[22]), .B(A[22]), .Z(n123) );
  COR2XL U109 ( .A(B[18]), .B(A[18]), .Z(n150) );
  COR2XL U110 ( .A(B[23]), .B(A[23]), .Z(n116) );
  CANR1XL U111 ( .A(n63), .B(n1), .C(n58), .Z(n61) );
  CENXL U112 ( .A(n61), .B(n62), .Z(SUM[30]) );
  COR2XL U113 ( .A(B[24]), .B(A[24]), .Z(n107) );
  COR2XL U114 ( .A(B[1]), .B(A[1]), .Z(n143) );
  COR2XL U115 ( .A(B[19]), .B(A[19]), .Z(n139) );
  COR2XL U116 ( .A(B[16]), .B(A[16]), .Z(n156) );
  COR2XL U117 ( .A(B[25]), .B(A[25]), .Z(n92) );
  CND2XL U118 ( .A(n78), .B(n79), .Z(n77) );
  COR2XL U119 ( .A(B[29]), .B(A[29]), .Z(n66) );
  COR2XL U120 ( .A(B[28]), .B(A[28]), .Z(n78) );
  COR2XL U121 ( .A(B[30]), .B(A[30]), .Z(n59) );
  CEOXL U122 ( .A(n46), .B(n47), .Z(SUM[3]) );
  COR2XL U123 ( .A(B[4]), .B(A[4]), .Z(n44) );
  CANR1XL U124 ( .A(n26), .B(n27), .C(n28), .Z(n23) );
  CNR2X1 U125 ( .A(n4), .B(n164), .Z(n163) );
  CND2X1 U126 ( .A(n208), .B(n209), .Z(n176) );
  CNR2X1 U127 ( .A(n210), .B(n199), .Z(n209) );
  CNR2X1 U128 ( .A(n212), .B(n213), .Z(n208) );
  CNR2IX1 U129 ( .B(n231), .A(n238), .Z(n236) );
  CNR2IX1 U130 ( .B(n239), .A(n240), .Z(n238) );
  CANR1XL U131 ( .A(n26), .B(n27), .C(n28), .Z(n240) );
  CNR2XL U132 ( .A(n225), .B(n212), .Z(n227) );
  CNR2XL U133 ( .A(n177), .B(n213), .Z(n237) );
  CND2X1 U134 ( .A(n136), .B(n99), .Z(n111) );
  CNR2IXL U135 ( .B(n177), .A(n176), .Z(n165) );
  CNR2XL U136 ( .A(n178), .B(n179), .Z(n204) );
  CNR2XL U137 ( .A(n178), .B(n179), .Z(n206) );
  CNR2XL U138 ( .A(n176), .B(n192), .Z(n190) );
  CENX1 U139 ( .A(n16), .B(n17), .Z(SUM[9]) );
  CENX1 U140 ( .A(n161), .B(n104), .Z(SUM[16]) );
  CENX1 U141 ( .A(n236), .B(n237), .Z(SUM[12]) );
  COND3X1 U142 ( .A(n98), .B(n99), .C(n100), .D(n101), .Z(n56) );
  CNR2IX1 U143 ( .B(n106), .A(n5), .Z(n100) );
  COND1XL U144 ( .A(n137), .B(n138), .C(n139), .Z(n99) );
  COND1XL U145 ( .A(n69), .B(n70), .C(n71), .Z(n50) );
  CANR1XL U146 ( .A(n156), .B(n104), .C(n159), .Z(n157) );
  CND2X1 U147 ( .A(n139), .B(n140), .Z(n145) );
  CANR1XL U148 ( .A(n10), .B(n104), .C(n138), .Z(n144) );
  CND2X1 U149 ( .A(n150), .B(n148), .Z(n152) );
  CANR1XL U150 ( .A(n8), .B(n104), .C(n149), .Z(n151) );
  CANR1XL U151 ( .A(n50), .B(n51), .C(n52), .Z(n46) );
  CANR1XL U152 ( .A(n13), .B(n1), .C(n67), .Z(n74) );
  CENX1 U153 ( .A(n68), .B(n50), .Z(SUM[2]) );
  COND1XL U154 ( .A(n126), .B(n127), .C(n128), .Z(n122) );
  COND1XL U155 ( .A(n18), .B(n19), .C(n20), .Z(n17) );
  COND4CX1 U156 ( .A(n19), .B(n20), .C(n252), .D(n22), .Z(n250) );
  CENX1 U157 ( .A(n141), .B(n72), .Z(SUM[1]) );
  CND2X1 U158 ( .A(n143), .B(n71), .Z(n141) );
  CENX1 U159 ( .A(n87), .B(n88), .Z(SUM[27]) );
  CANR1XL U160 ( .A(n11), .B(n56), .C(n85), .Z(n87) );
  CNR2X1 U161 ( .A(n260), .B(n261), .Z(n241) );
  CNR2IX1 U162 ( .B(n20), .A(n18), .Z(n24) );
  CND2X1 U163 ( .A(n254), .B(n255), .Z(n28) );
  CND3XL U164 ( .A(n39), .B(n184), .C(n185), .Z(n255) );
  CENX1 U165 ( .A(n251), .B(n250), .Z(SUM[10]) );
  CENX1 U166 ( .A(n214), .B(n215), .Z(SUM[15]) );
  CNR2IXL U167 ( .B(n197), .A(n210), .Z(n215) );
  CANR1XL U168 ( .A(n217), .B(n218), .C(n219), .Z(n216) );
  CANR1XL U169 ( .A(n230), .B(n231), .C(n232), .Z(n229) );
  CND2X1 U170 ( .A(n235), .B(n231), .Z(n228) );
  CNR2IX1 U171 ( .B(n91), .A(n89), .Z(n95) );
  CANR1XL U172 ( .A(n92), .B(n56), .C(n96), .Z(n94) );
  CENX1 U173 ( .A(n131), .B(n132), .Z(SUM[21]) );
  CND2X1 U174 ( .A(n129), .B(n128), .Z(n131) );
  COND1XL U175 ( .A(n133), .B(n134), .C(n127), .Z(n132) );
  CND2X1 U176 ( .A(n142), .B(n71), .Z(n262) );
  CNR2X1 U177 ( .A(n264), .B(n69), .Z(n263) );
  CANR1XL U178 ( .A(n9), .B(n111), .C(n122), .Z(n124) );
  CND2X1 U179 ( .A(n107), .B(n106), .Z(n110) );
  CANR1XL U180 ( .A(n7), .B(n111), .C(n108), .Z(n109) );
  CND2X1 U181 ( .A(n116), .B(n114), .Z(n118) );
  CANR1XL U182 ( .A(n6), .B(n111), .C(n115), .Z(n117) );
  CEOXL U183 ( .A(n3), .B(n41), .Z(SUM[5]) );
  CND2X1 U184 ( .A(n39), .B(n38), .Z(n41) );
  CANR1XL U185 ( .A(n33), .B(n34), .C(n35), .Z(n29) );
  CND2X1 U186 ( .A(n20), .B(n22), .Z(n172) );
  CENX1 U187 ( .A(n226), .B(n227), .Z(SUM[13]) );
  CNR2XL U188 ( .A(n199), .B(n200), .Z(n195) );
  CND2X1 U189 ( .A(n7), .B(n107), .Z(n98) );
  CNR2IX1 U190 ( .B(n59), .A(n60), .Z(n55) );
  CNR2XL U191 ( .A(n176), .B(n179), .Z(n180) );
  CND3XL U192 ( .A(n39), .B(n184), .C(n185), .Z(n183) );
  CND3XL U193 ( .A(n21), .B(n25), .C(n234), .Z(n230) );
  CND2X1 U194 ( .A(n52), .B(n49), .Z(n192) );
  CND2X1 U195 ( .A(n156), .B(n160), .Z(n161) );
  CAN2X1 U196 ( .A(n9), .B(n123), .Z(n6) );
  CAN2X1 U197 ( .A(n6), .B(n116), .Z(n7) );
  CAN2X1 U198 ( .A(n156), .B(n155), .Z(n8) );
  CAN2X1 U199 ( .A(n130), .B(n129), .Z(n9) );
  CAN2X1 U200 ( .A(n8), .B(n150), .Z(n10) );
  CAN2X1 U201 ( .A(n92), .B(n93), .Z(n11) );
  CAN2X1 U202 ( .A(n11), .B(n86), .Z(n12) );
  CAN2X1 U203 ( .A(n12), .B(n78), .Z(n13) );
  CAN2X1 U204 ( .A(n35), .B(n31), .Z(n14) );
  CND2X1 U205 ( .A(n13), .B(n66), .Z(n60) );
  CNR2IX1 U206 ( .B(n32), .A(n14), .Z(n182) );
  CND2X1 U207 ( .A(n174), .B(n249), .Z(n247) );
  CND2X1 U208 ( .A(n10), .B(n139), .Z(n105) );
  CND2X1 U209 ( .A(n220), .B(n211), .Z(n219) );
  CNR2X1 U210 ( .A(n243), .B(n244), .Z(n242) );
  CND2X1 U211 ( .A(n21), .B(n25), .Z(n243) );
  CND2X1 U212 ( .A(n197), .B(n198), .Z(n196) );
  CNR2X1 U213 ( .A(n258), .B(n259), .Z(n257) );
  CND2X1 U214 ( .A(n34), .B(n31), .Z(n259) );
  COND1XL U215 ( .A(n82), .B(n83), .C(n84), .Z(n79) );
  CND2X1 U216 ( .A(n171), .B(n172), .Z(n170) );
  CND2XL U217 ( .A(n34), .B(n40), .Z(n36) );
  COND2XL U218 ( .A(A[10]), .B(B[10]), .C(A[9]), .D(B[9]), .Z(n246) );
  CEOXL U219 ( .A(B[29]), .B(A[29]), .Z(n75) );
  CENX1 U220 ( .A(n80), .B(n81), .Z(SUM[28]) );
  CEOXL U221 ( .A(B[28]), .B(A[28]), .Z(n81) );
  CANR1XL U222 ( .A(n12), .B(n1), .C(n79), .Z(n80) );
  CAOR1X1 U223 ( .A(n59), .B(n58), .C(n15), .Z(n57) );
  CAN2XL U224 ( .A(B[30]), .B(A[30]), .Z(n15) );
  CND2XL U225 ( .A(B[20]), .B(A[20]), .Z(n127) );
  CND2XL U226 ( .A(B[11]), .B(A[11]), .Z(n173) );
  CND2XL U227 ( .A(B[25]), .B(A[25]), .Z(n90) );
  CND2XL U228 ( .A(B[13]), .B(A[13]), .Z(n200) );
  CND2XL U229 ( .A(B[23]), .B(A[23]), .Z(n114) );
  CND2XL U230 ( .A(B[18]), .B(A[18]), .Z(n148) );
  CND2XL U231 ( .A(B[17]), .B(A[17]), .Z(n153) );
  CND2X1 U232 ( .A(n64), .B(n65), .Z(n58) );
  CND2XL U233 ( .A(B[29]), .B(A[29]), .Z(n64) );
  CND2X1 U234 ( .A(n66), .B(n67), .Z(n65) );
  CND2X1 U235 ( .A(n153), .B(n154), .Z(n149) );
  CND3XL U236 ( .A(A[16]), .B(B[16]), .C(n155), .Z(n154) );
  CND2XL U237 ( .A(B[19]), .B(A[19]), .Z(n140) );
  CND2XL U238 ( .A(B[16]), .B(A[16]), .Z(n160) );
  CND2XL U239 ( .A(B[26]), .B(A[26]), .Z(n91) );
  CND2XL U240 ( .A(B[27]), .B(A[27]), .Z(n84) );
  CND2XL U241 ( .A(B[24]), .B(A[24]), .Z(n106) );
  CANR1X1 U242 ( .A(n55), .B(n56), .C(n57), .Z(n53) );
  CND2X1 U243 ( .A(n76), .B(n77), .Z(n67) );
  CND2X1 U244 ( .A(n266), .B(n267), .Z(n265) );
  CENX1 U245 ( .A(n45), .B(n27), .Z(SUM[4]) );
  CENX1 U246 ( .A(n23), .B(n24), .Z(SUM[8]) );
  CEOXL U247 ( .A(B[30]), .B(A[30]), .Z(n62) );
  CIVX2 U248 ( .A(n142), .Z(n72) );
  CIVX2 U249 ( .A(n48), .Z(n260) );
  CND2XL U250 ( .A(B[28]), .B(A[28]), .Z(n76) );
  COND2XL U251 ( .A(A[7]), .B(B[7]), .C(A[6]), .D(B[6]), .Z(n256) );
  CEOXL U252 ( .A(B[31]), .B(A[31]), .Z(n54) );
  CND2XL U253 ( .A(B[22]), .B(A[22]), .Z(n121) );
  CND2X1 U254 ( .A(n123), .B(n121), .Z(n125) );
  CIVX2 U255 ( .A(n39), .Z(n37) );
  CIVX2 U256 ( .A(n60), .Z(n63) );
  CIVX2 U257 ( .A(n72), .Z(n70) );
  CIVX2 U258 ( .A(n85), .Z(n83) );
  CIVX2 U259 ( .A(n86), .Z(n82) );
  CIVX2 U260 ( .A(n93), .Z(n89) );
  CIVX2 U261 ( .A(n90), .Z(n96) );
  CIVX2 U262 ( .A(n105), .Z(n103) );
  CIVX2 U263 ( .A(n98), .Z(n102) );
  CIVX2 U264 ( .A(n116), .Z(n112) );
  CIVX2 U265 ( .A(n123), .Z(n119) );
  CIVX2 U266 ( .A(n129), .Z(n126) );
  CIVX2 U267 ( .A(n130), .Z(n133) );
  CIVX2 U268 ( .A(n111), .Z(n134) );
  CIVX2 U269 ( .A(n140), .Z(n137) );
  CND2IX1 U270 ( .B(n105), .A(n104), .Z(n136) );
  CIVX2 U271 ( .A(n150), .Z(n146) );
  CIVX2 U272 ( .A(n160), .Z(n159) );
  CND2IX1 U273 ( .B(n165), .A(n166), .Z(n164) );
  CND2X1 U274 ( .A(n167), .B(n168), .Z(n166) );
  CND2IX1 U275 ( .B(n169), .A(n170), .Z(n168) );
  CND2X1 U276 ( .A(n182), .B(n183), .Z(n181) );
  CND2IX1 U277 ( .B(n188), .A(n189), .Z(n187) );
  CND2X1 U278 ( .A(n190), .B(n191), .Z(n189) );
  CND2X1 U279 ( .A(n201), .B(n202), .Z(n186) );
  CND2X1 U280 ( .A(n205), .B(n206), .Z(n201) );
  CIVX2 U281 ( .A(n211), .Z(n199) );
  CIVX2 U282 ( .A(n193), .Z(n210) );
  CAN2X1 U283 ( .A(n221), .B(n200), .Z(n217) );
  CIVX2 U284 ( .A(n220), .Z(n212) );
  CIVX2 U285 ( .A(n200), .Z(n225) );
  CIVX2 U286 ( .A(n28), .Z(n235) );
  CIVX2 U287 ( .A(n233), .Z(n213) );
  CIVX2 U288 ( .A(n221), .Z(n177) );
  CIVX2 U289 ( .A(n241), .Z(n27) );
  CIVX2 U290 ( .A(n178), .Z(n26) );
  CIVX2 U291 ( .A(n179), .Z(n239) );
  CIVX2 U292 ( .A(n242), .Z(n179) );
  CIVX2 U293 ( .A(n256), .Z(n184) );
  CIVX2 U294 ( .A(n40), .Z(n35) );
  CIVX2 U295 ( .A(n257), .Z(n178) );
  CIVX2 U296 ( .A(n73), .Z(n52) );
  CIVX2 U297 ( .A(n143), .Z(n69) );
  CIVX2 U298 ( .A(n51), .Z(n264) );
  CIVX2 U299 ( .A(A[0]), .Z(n267) );
endmodule


module nios_2_DW01_add_6 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265;

  CND2XL U2 ( .A(n40), .B(n39), .Z(n42) );
  CIVX1 U3 ( .A(n40), .Z(n38) );
  CENXL U4 ( .A(n74), .B(n75), .Z(SUM[29]) );
  COND3X1 U5 ( .A(n98), .B(n99), .C(n100), .D(n101), .Z(n56) );
  CND3X1 U6 ( .A(n102), .B(n103), .C(n104), .Z(n101) );
  COND1XL U7 ( .A(n120), .B(n121), .C(n122), .Z(n116) );
  CANR1X1 U8 ( .A(n55), .B(n56), .C(n57), .Z(n53) );
  CND2X1 U9 ( .A(n175), .B(n247), .Z(n245) );
  CAN2XL U10 ( .A(n263), .B(n143), .Z(SUM[0]) );
  CEOXL U11 ( .A(n30), .B(n31), .Z(SUM[7]) );
  CENXL U12 ( .A(n97), .B(n56), .Z(SUM[25]) );
  CENXL U13 ( .A(n53), .B(n54), .Z(SUM[31]) );
  CND2XL U14 ( .A(n22), .B(n26), .Z(n250) );
  COR2X1 U15 ( .A(B[8]), .B(A[8]), .Z(n26) );
  COR2XL U16 ( .A(B[18]), .B(A[18]), .Z(n151) );
  COR2X1 U17 ( .A(B[17]), .B(A[17]), .Z(n156) );
  COR2XL U18 ( .A(B[15]), .B(A[15]), .Z(n192) );
  CAN2XL U19 ( .A(n92), .B(n93), .Z(n11) );
  CNR2IXL U20 ( .B(n176), .A(n177), .Z(n168) );
  COND1XL U21 ( .A(n147), .B(n148), .C(n149), .Z(n139) );
  CNR2X1 U22 ( .A(n5), .B(n165), .Z(n164) );
  CNR2XL U23 ( .A(n179), .B(n180), .Z(n190) );
  CNR2XL U24 ( .A(n177), .B(n206), .Z(n204) );
  CAN2XL U25 ( .A(n2), .B(n3), .Z(n5) );
  CND2XL U26 ( .A(n181), .B(n182), .Z(n3) );
  COND1XL U27 ( .A(n138), .B(n139), .C(n140), .Z(n99) );
  CENX1 U28 ( .A(n245), .B(n246), .Z(SUM[11]) );
  CNR2IX1 U29 ( .B(n197), .A(n215), .Z(n213) );
  CEOXL U30 ( .A(n152), .B(n153), .Z(SUM[18]) );
  CNR2XL U31 ( .A(n251), .B(n29), .Z(n20) );
  CNR2XL U32 ( .A(n177), .B(n180), .Z(n2) );
  CND2X2 U33 ( .A(n163), .B(n164), .Z(n104) );
  CNR2XL U34 ( .A(n179), .B(n180), .Z(n205) );
  CND2XL U35 ( .A(n32), .B(n33), .Z(n31) );
  COND4CXL U36 ( .A(n172), .B(n173), .C(n243), .D(n176), .Z(n230) );
  CND2XL U37 ( .A(n174), .B(n175), .Z(n243) );
  CND2X2 U38 ( .A(n7), .B(n108), .Z(n98) );
  CND2XL U39 ( .A(n206), .B(n191), .Z(n259) );
  CNR2XL U40 ( .A(n258), .B(n259), .Z(n239) );
  CEOXL U41 ( .A(n125), .B(n126), .Z(SUM[22]) );
  CEOXL U42 ( .A(n118), .B(n119), .Z(SUM[23]) );
  CNR2IXL U43 ( .B(n84), .A(n82), .Z(n88) );
  CNR2IXL U44 ( .B(n91), .A(n89), .Z(n95) );
  CNR2IXL U45 ( .B(n33), .A(n14), .Z(n252) );
  CND2XL U46 ( .A(n131), .B(n128), .Z(n136) );
  CAN2X1 U47 ( .A(n43), .B(n4), .Z(n15) );
  CND2X1 U48 ( .A(n44), .B(n28), .Z(n4) );
  CND2XL U49 ( .A(n92), .B(n90), .Z(n97) );
  CND2XL U50 ( .A(n130), .B(n129), .Z(n132) );
  CND2XL U51 ( .A(n233), .B(n175), .Z(n249) );
  CND2XL U52 ( .A(n51), .B(n73), .Z(n68) );
  CND2XL U53 ( .A(n144), .B(n71), .Z(n142) );
  CND2XL U54 ( .A(n140), .B(n141), .Z(n146) );
  CND2XL U55 ( .A(n151), .B(n149), .Z(n153) );
  CNR2XL U56 ( .A(n48), .B(n177), .Z(n202) );
  CNR2XL U57 ( .A(n179), .B(n180), .Z(n203) );
  CND2XL U58 ( .A(n196), .B(n197), .Z(n195) );
  CND2XL U59 ( .A(n174), .B(n176), .Z(n246) );
  CEOXL U60 ( .A(n221), .B(n222), .Z(SUM[14]) );
  CND2XL U61 ( .A(n210), .B(n197), .Z(n222) );
  CEOXL U62 ( .A(n110), .B(n111), .Z(SUM[24]) );
  CND2XL U63 ( .A(n48), .B(n49), .Z(n47) );
  CND2XL U64 ( .A(n156), .B(n154), .Z(n159) );
  CIVXL U65 ( .A(n150), .Z(n148) );
  CIVXL U66 ( .A(n123), .Z(n121) );
  COND1X1 U67 ( .A(n113), .B(n114), .C(n115), .Z(n109) );
  CIVXL U68 ( .A(n116), .Z(n114) );
  COR2XL U69 ( .A(B[11]), .B(A[11]), .Z(n176) );
  COR2XL U70 ( .A(B[5]), .B(A[5]), .Z(n40) );
  CND2XL U71 ( .A(B[9]), .B(A[9]), .Z(n23) );
  CND2XL U72 ( .A(B[8]), .B(A[8]), .Z(n21) );
  COR2XL U73 ( .A(B[14]), .B(A[14]), .Z(n210) );
  COR2XL U74 ( .A(B[13]), .B(A[13]), .Z(n219) );
  CND2XL U75 ( .A(B[5]), .B(A[5]), .Z(n39) );
  COR2XL U76 ( .A(B[21]), .B(A[21]), .Z(n130) );
  COR2XL U77 ( .A(B[22]), .B(A[22]), .Z(n124) );
  COR2XL U78 ( .A(B[23]), .B(A[23]), .Z(n117) );
  COR2XL U79 ( .A(B[20]), .B(A[20]), .Z(n131) );
  COR2XL U80 ( .A(B[10]), .B(A[10]), .Z(n233) );
  COR2XL U81 ( .A(B[9]), .B(A[9]), .Z(n22) );
  COR2XL U82 ( .A(B[24]), .B(A[24]), .Z(n108) );
  COR2XL U83 ( .A(B[12]), .B(A[12]), .Z(n232) );
  COR2XL U84 ( .A(B[7]), .B(A[7]), .Z(n32) );
  COR2XL U85 ( .A(B[4]), .B(A[4]), .Z(n44) );
  COR2XL U86 ( .A(B[1]), .B(A[1]), .Z(n144) );
  COR2XL U87 ( .A(B[26]), .B(A[26]), .Z(n93) );
  COR2XL U88 ( .A(B[27]), .B(A[27]), .Z(n86) );
  COR2XL U89 ( .A(B[3]), .B(A[3]), .Z(n49) );
  COR2XL U90 ( .A(B[19]), .B(A[19]), .Z(n140) );
  COR2XL U91 ( .A(B[16]), .B(A[16]), .Z(n157) );
  COR2XL U92 ( .A(B[25]), .B(A[25]), .Z(n92) );
  CND2XL U93 ( .A(n78), .B(n79), .Z(n77) );
  COR2XL U94 ( .A(B[29]), .B(A[29]), .Z(n66) );
  COR2XL U95 ( .A(B[28]), .B(A[28]), .Z(n78) );
  COR2XL U96 ( .A(B[6]), .B(A[6]), .Z(n35) );
  COR2XL U97 ( .A(B[30]), .B(A[30]), .Z(n59) );
  CND2XL U98 ( .A(B[4]), .B(A[4]), .Z(n43) );
  CNR2XL U99 ( .A(n239), .B(n179), .Z(n251) );
  CANR1XL U100 ( .A(n10), .B(n104), .C(n139), .Z(n145) );
  CANR1XL U101 ( .A(n11), .B(n56), .C(n85), .Z(n87) );
  CANR1XL U102 ( .A(n12), .B(n56), .C(n79), .Z(n80) );
  CENX1 U103 ( .A(n94), .B(n95), .Z(SUM[26]) );
  CNR2X1 U104 ( .A(n185), .B(n186), .Z(n163) );
  CND2X1 U105 ( .A(n207), .B(n208), .Z(n177) );
  CNR2X1 U106 ( .A(n209), .B(n198), .Z(n208) );
  CNR2X1 U107 ( .A(n211), .B(n212), .Z(n207) );
  CENX1 U108 ( .A(n87), .B(n88), .Z(SUM[27]) );
  CANR1XL U109 ( .A(n27), .B(n28), .C(n29), .Z(n238) );
  CENX1 U110 ( .A(n235), .B(n236), .Z(SUM[12]) );
  CNR2XL U111 ( .A(n178), .B(n212), .Z(n236) );
  CNR2IX1 U112 ( .B(n230), .A(n237), .Z(n235) );
  CNR2IX1 U113 ( .B(n240), .A(n238), .Z(n237) );
  CND2X1 U114 ( .A(n137), .B(n99), .Z(n112) );
  CNR2IXL U115 ( .B(n178), .A(n177), .Z(n166) );
  CENX1 U116 ( .A(n132), .B(n133), .Z(SUM[21]) );
  CNR2XL U117 ( .A(n177), .B(n191), .Z(n189) );
  CENX1 U118 ( .A(n249), .B(n248), .Z(SUM[10]) );
  CEOX1 U119 ( .A(n145), .B(n146), .Z(SUM[19]) );
  CAN2X1 U120 ( .A(n106), .B(n107), .Z(n100) );
  COND1XL U121 ( .A(n38), .B(n15), .C(n39), .Z(n34) );
  COND1XL U122 ( .A(n69), .B(n70), .C(n71), .Z(n50) );
  CANR1XL U123 ( .A(n9), .B(n104), .C(n150), .Z(n152) );
  CEOX1 U124 ( .A(n46), .B(n47), .Z(SUM[3]) );
  CANR1XL U125 ( .A(n50), .B(n51), .C(n52), .Z(n46) );
  CANR1XL U126 ( .A(n63), .B(n56), .C(n58), .Z(n61) );
  CANR1XL U127 ( .A(n92), .B(n56), .C(n96), .Z(n94) );
  COND1X1 U128 ( .A(n89), .B(n90), .C(n91), .Z(n85) );
  COND1XL U129 ( .A(n127), .B(n128), .C(n129), .Z(n123) );
  COND1XL U130 ( .A(n134), .B(n135), .C(n128), .Z(n133) );
  COND4CX1 U131 ( .A(n20), .B(n21), .C(n250), .D(n23), .Z(n248) );
  CENXL U132 ( .A(n61), .B(n62), .Z(SUM[30]) );
  CENX1 U133 ( .A(n80), .B(n81), .Z(SUM[28]) );
  CENX1 U134 ( .A(n37), .B(n34), .Z(SUM[6]) );
  CND2XL U135 ( .A(n35), .B(n41), .Z(n37) );
  CENX1 U136 ( .A(n162), .B(n104), .Z(SUM[16]) );
  CND2X1 U137 ( .A(n157), .B(n161), .Z(n162) );
  CENX1 U138 ( .A(n17), .B(n18), .Z(SUM[9]) );
  CND2X1 U139 ( .A(n22), .B(n23), .Z(n17) );
  COND1XL U140 ( .A(n19), .B(n20), .C(n21), .Z(n18) );
  CANR1XL U141 ( .A(n216), .B(n217), .C(n218), .Z(n215) );
  CND2X1 U142 ( .A(n219), .B(n210), .Z(n218) );
  CEOX1 U143 ( .A(n135), .B(n136), .Z(SUM[20]) );
  CND2X1 U144 ( .A(n252), .B(n253), .Z(n29) );
  CND3XL U145 ( .A(n40), .B(n183), .C(n184), .Z(n253) );
  CANR1XL U146 ( .A(n34), .B(n35), .C(n36), .Z(n30) );
  COND4CX1 U147 ( .A(n27), .B(n28), .C(n227), .D(n228), .Z(n217) );
  CANR1XL U148 ( .A(n229), .B(n230), .C(n231), .Z(n228) );
  CND2X1 U149 ( .A(n234), .B(n230), .Z(n227) );
  CND2X1 U150 ( .A(n176), .B(n232), .Z(n231) );
  CND3XL U151 ( .A(n49), .B(n260), .C(n261), .Z(n206) );
  CND2X1 U152 ( .A(n143), .B(n71), .Z(n260) );
  CNR2X1 U153 ( .A(n262), .B(n69), .Z(n261) );
  CANR1XL U154 ( .A(n8), .B(n112), .C(n123), .Z(n125) );
  CND2X1 U155 ( .A(n117), .B(n115), .Z(n119) );
  CANR1XL U156 ( .A(n6), .B(n112), .C(n116), .Z(n118) );
  CND2X1 U157 ( .A(n21), .B(n23), .Z(n173) );
  CNR2XL U158 ( .A(n198), .B(n199), .Z(n194) );
  CENX1 U159 ( .A(n68), .B(n50), .Z(SUM[2]) );
  CNR2IX1 U160 ( .B(n59), .A(n60), .Z(n55) );
  CND2X1 U161 ( .A(n108), .B(n106), .Z(n111) );
  CANR1XL U162 ( .A(n7), .B(n112), .C(n109), .Z(n110) );
  CNR2IX1 U163 ( .B(n192), .A(n193), .Z(n187) );
  CNR2X1 U164 ( .A(n194), .B(n195), .Z(n193) );
  CND3XL U165 ( .A(n22), .B(n26), .C(n233), .Z(n229) );
  CND2X1 U166 ( .A(n43), .B(n39), .Z(n184) );
  CENX1 U167 ( .A(n142), .B(n72), .Z(SUM[1]) );
  CND2X1 U168 ( .A(n52), .B(n49), .Z(n191) );
  CND3XL U169 ( .A(n40), .B(n183), .C(n184), .Z(n182) );
  CAN2X1 U170 ( .A(n8), .B(n124), .Z(n6) );
  CAN2X1 U171 ( .A(n6), .B(n117), .Z(n7) );
  CAN2X1 U172 ( .A(n131), .B(n130), .Z(n8) );
  CAN2X1 U173 ( .A(n157), .B(n156), .Z(n9) );
  CAN2X1 U174 ( .A(n9), .B(n151), .Z(n10) );
  CAN2X1 U175 ( .A(n11), .B(n86), .Z(n12) );
  CAN2X1 U176 ( .A(n12), .B(n78), .Z(n13) );
  CAN2X1 U177 ( .A(n36), .B(n32), .Z(n14) );
  CND2X1 U178 ( .A(n13), .B(n66), .Z(n60) );
  CNR2IX1 U179 ( .B(n33), .A(n14), .Z(n181) );
  CND2X1 U180 ( .A(n10), .B(n140), .Z(n105) );
  CND2X1 U181 ( .A(n233), .B(n248), .Z(n247) );
  CNR2X1 U182 ( .A(n241), .B(n242), .Z(n240) );
  CND2X1 U183 ( .A(n22), .B(n26), .Z(n241) );
  CND2X1 U184 ( .A(n176), .B(n233), .Z(n242) );
  CNR2X1 U185 ( .A(n256), .B(n257), .Z(n255) );
  CND2X1 U186 ( .A(n35), .B(n32), .Z(n257) );
  CND2X1 U187 ( .A(n40), .B(n44), .Z(n256) );
  CND2X1 U188 ( .A(n108), .B(n109), .Z(n107) );
  CEOX1 U189 ( .A(n158), .B(n159), .Z(SUM[17]) );
  CANR1XL U190 ( .A(n157), .B(n104), .C(n160), .Z(n158) );
  CENX1 U191 ( .A(n225), .B(n226), .Z(SUM[13]) );
  CNR2XL U192 ( .A(n224), .B(n211), .Z(n226) );
  CNR2IX1 U193 ( .B(n220), .A(n223), .Z(n225) );
  COND1XL U194 ( .A(n82), .B(n83), .C(n84), .Z(n79) );
  CND2X1 U195 ( .A(n172), .B(n173), .Z(n171) );
  CANR4CX1 U196 ( .A(n178), .B(n223), .C(n219), .D(n224), .Z(n221) );
  CND2X1 U197 ( .A(n174), .B(n175), .Z(n170) );
  CENX1 U198 ( .A(n213), .B(n214), .Z(SUM[15]) );
  CNR2IXL U199 ( .B(n196), .A(n209), .Z(n214) );
  CEOXL U200 ( .A(n15), .B(n42), .Z(SUM[5]) );
  CENX1 U201 ( .A(n45), .B(n28), .Z(SUM[4]) );
  CND2X1 U202 ( .A(n44), .B(n43), .Z(n45) );
  CENX1 U203 ( .A(n24), .B(n25), .Z(SUM[8]) );
  CNR2IX1 U204 ( .B(n21), .A(n19), .Z(n25) );
  CANR1XL U205 ( .A(n27), .B(n28), .C(n29), .Z(n24) );
  COND2XL U206 ( .A(A[10]), .B(B[10]), .C(A[9]), .D(B[9]), .Z(n244) );
  CEOXL U207 ( .A(B[28]), .B(A[28]), .Z(n81) );
  CEOXL U208 ( .A(B[29]), .B(A[29]), .Z(n75) );
  CANR1XL U209 ( .A(n13), .B(n56), .C(n67), .Z(n74) );
  CND2XL U210 ( .A(B[10]), .B(A[10]), .Z(n175) );
  CAOR1X1 U211 ( .A(n59), .B(n58), .C(n16), .Z(n57) );
  CAN2XL U212 ( .A(B[30]), .B(A[30]), .Z(n16) );
  CND2XL U213 ( .A(B[1]), .B(A[1]), .Z(n71) );
  CND2XL U214 ( .A(B[20]), .B(A[20]), .Z(n128) );
  CND2XL U215 ( .A(B[0]), .B(A[0]), .Z(n143) );
  CND2XL U216 ( .A(B[11]), .B(A[11]), .Z(n174) );
  CND2XL U217 ( .A(B[25]), .B(A[25]), .Z(n90) );
  CND2XL U218 ( .A(B[3]), .B(A[3]), .Z(n48) );
  CND2XL U219 ( .A(B[14]), .B(A[14]), .Z(n197) );
  CND2XL U220 ( .A(B[13]), .B(A[13]), .Z(n199) );
  CND2XL U221 ( .A(B[21]), .B(A[21]), .Z(n129) );
  CND2XL U222 ( .A(B[18]), .B(A[18]), .Z(n149) );
  CND2XL U223 ( .A(B[23]), .B(A[23]), .Z(n115) );
  CND2XL U224 ( .A(B[17]), .B(A[17]), .Z(n154) );
  CND2X1 U225 ( .A(n64), .B(n65), .Z(n58) );
  CND2XL U226 ( .A(B[29]), .B(A[29]), .Z(n64) );
  CND2X1 U227 ( .A(n66), .B(n67), .Z(n65) );
  CND2X1 U228 ( .A(n154), .B(n155), .Z(n150) );
  CND3XL U229 ( .A(A[16]), .B(B[16]), .C(n156), .Z(n155) );
  CND2XL U230 ( .A(B[7]), .B(A[7]), .Z(n33) );
  CND2XL U231 ( .A(B[2]), .B(A[2]), .Z(n73) );
  CND2XL U232 ( .A(B[19]), .B(A[19]), .Z(n141) );
  CND2XL U233 ( .A(B[16]), .B(A[16]), .Z(n161) );
  CND2XL U234 ( .A(B[12]), .B(A[12]), .Z(n220) );
  CND2XL U235 ( .A(B[26]), .B(A[26]), .Z(n91) );
  CND2XL U236 ( .A(B[27]), .B(A[27]), .Z(n84) );
  CND2XL U237 ( .A(B[24]), .B(A[24]), .Z(n106) );
  CND2XL U238 ( .A(B[15]), .B(A[15]), .Z(n196) );
  CND2X1 U239 ( .A(n76), .B(n77), .Z(n67) );
  CND2X1 U240 ( .A(n264), .B(n265), .Z(n263) );
  COR2X1 U241 ( .A(B[2]), .B(A[2]), .Z(n51) );
  CEOXL U242 ( .A(B[30]), .B(A[30]), .Z(n62) );
  CIVX2 U243 ( .A(n143), .Z(n72) );
  CIVX2 U244 ( .A(n48), .Z(n258) );
  CND2XL U245 ( .A(B[28]), .B(A[28]), .Z(n76) );
  COND2XL U246 ( .A(A[7]), .B(B[7]), .C(A[6]), .D(B[6]), .Z(n254) );
  CND2XL U247 ( .A(B[6]), .B(A[6]), .Z(n41) );
  CEOXL U248 ( .A(B[31]), .B(A[31]), .Z(n54) );
  CND2X1 U249 ( .A(B[22]), .B(A[22]), .Z(n122) );
  CND2X1 U250 ( .A(n124), .B(n122), .Z(n126) );
  CIVX2 U251 ( .A(n26), .Z(n19) );
  CIVX2 U252 ( .A(n60), .Z(n63) );
  CIVX2 U253 ( .A(n72), .Z(n70) );
  CIVX2 U254 ( .A(n85), .Z(n83) );
  CIVX2 U255 ( .A(n86), .Z(n82) );
  CIVX2 U256 ( .A(n93), .Z(n89) );
  CIVX2 U257 ( .A(n90), .Z(n96) );
  CIVX2 U258 ( .A(n105), .Z(n103) );
  CIVX2 U259 ( .A(n98), .Z(n102) );
  CIVX2 U260 ( .A(n117), .Z(n113) );
  CIVX2 U261 ( .A(n124), .Z(n120) );
  CIVX2 U262 ( .A(n130), .Z(n127) );
  CIVX2 U263 ( .A(n131), .Z(n134) );
  CIVX2 U264 ( .A(n112), .Z(n135) );
  CIVX2 U265 ( .A(n141), .Z(n138) );
  CND2IX1 U266 ( .B(n105), .A(n104), .Z(n137) );
  CIVX2 U267 ( .A(n151), .Z(n147) );
  CIVX2 U268 ( .A(n161), .Z(n160) );
  CND2IX1 U269 ( .B(n166), .A(n167), .Z(n165) );
  CND2X1 U270 ( .A(n168), .B(n169), .Z(n167) );
  CND2IX1 U271 ( .B(n170), .A(n171), .Z(n169) );
  CND2IX1 U272 ( .B(n187), .A(n188), .Z(n186) );
  CND2X1 U273 ( .A(n189), .B(n190), .Z(n188) );
  CND2X1 U274 ( .A(n200), .B(n201), .Z(n185) );
  CND2X1 U275 ( .A(n202), .B(n203), .Z(n201) );
  CND2X1 U276 ( .A(n204), .B(n205), .Z(n200) );
  CIVX2 U277 ( .A(n210), .Z(n198) );
  CIVX2 U278 ( .A(n192), .Z(n209) );
  CAN2X1 U279 ( .A(n220), .B(n199), .Z(n216) );
  CIVX2 U280 ( .A(n219), .Z(n211) );
  CIVX2 U281 ( .A(n199), .Z(n224) );
  CIVX2 U282 ( .A(n217), .Z(n223) );
  CIVX2 U283 ( .A(n29), .Z(n234) );
  CIVX2 U284 ( .A(n232), .Z(n212) );
  CIVX2 U285 ( .A(n220), .Z(n178) );
  CIVX2 U286 ( .A(n239), .Z(n28) );
  CIVX2 U287 ( .A(n179), .Z(n27) );
  CIVX2 U288 ( .A(n240), .Z(n180) );
  CIVX2 U289 ( .A(n244), .Z(n172) );
  CIVX2 U290 ( .A(n254), .Z(n183) );
  CIVX2 U291 ( .A(n41), .Z(n36) );
  CIVX2 U292 ( .A(n255), .Z(n179) );
  CIVX2 U293 ( .A(n73), .Z(n52) );
  CIVX2 U294 ( .A(n144), .Z(n69) );
  CIVX2 U295 ( .A(n51), .Z(n262) );
  CIVX2 U296 ( .A(A[0]), .Z(n265) );
  CIVX2 U297 ( .A(B[0]), .Z(n264) );
endmodule


module nios_2_DW01_add_10 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160;

  CNR2X1 U2 ( .A(n139), .B(n140), .Z(n138) );
  CNR2X1 U3 ( .A(n130), .B(n131), .Z(n129) );
  CNIVX1 U4 ( .A(B[14]), .Z(n1) );
  CNIVX1 U5 ( .A(B[12]), .Z(n2) );
  CNIVX1 U6 ( .A(B[8]), .Z(n3) );
  CNIVX1 U7 ( .A(B[20]), .Z(n4) );
  CNIVX1 U8 ( .A(B[17]), .Z(n5) );
  CNIVXL U9 ( .A(B[13]), .Z(n6) );
  CNIVXL U10 ( .A(B[21]), .Z(n7) );
  CNIVX1 U11 ( .A(B[9]), .Z(n8) );
  CND3X1 U12 ( .A(n6), .B(n2), .C(n122), .Z(n9) );
  CNIVXL U13 ( .A(B[26]), .Z(n10) );
  CNIVXL U14 ( .A(B[18]), .Z(n11) );
  CNIVXL U15 ( .A(B[25]), .Z(n12) );
  CNIVXL U16 ( .A(B[15]), .Z(n13) );
  CNIVX1 U17 ( .A(B[16]), .Z(n14) );
  CENX1 U18 ( .A(n60), .B(n15), .Z(SUM[4]) );
  CEOX1 U19 ( .A(n13), .B(n18), .Z(SUM[15]) );
  CNR2X1 U20 ( .A(n121), .B(n9), .Z(n18) );
  COND1X1 U21 ( .A(n41), .B(n57), .C(n58), .Z(n54) );
  CNR2XL U22 ( .A(n99), .B(n100), .Z(n17) );
  CEOXL U23 ( .A(B[22]), .B(n17), .Z(SUM[22]) );
  CEOX1 U24 ( .A(n127), .B(n129), .Z(SUM[11]) );
  CAN2X2 U25 ( .A(n22), .B(n91), .Z(n72) );
  CAN2XL U26 ( .A(n24), .B(n91), .Z(n23) );
  CNR2XL U27 ( .A(A[2]), .B(B[2]), .Z(n146) );
  CIVXL U28 ( .A(B[27]), .Z(n90) );
  CND2XL U29 ( .A(n33), .B(n41), .Z(n126) );
  CND2XL U30 ( .A(n26), .B(n23), .Z(n93) );
  CND2XL U31 ( .A(n59), .B(n58), .Z(n15) );
  CAN2XL U32 ( .A(n25), .B(n4), .Z(n24) );
  CENX1 U33 ( .A(n16), .B(n4), .Z(SUM[20]) );
  CND2XL U34 ( .A(n25), .B(n91), .Z(n16) );
  CND2XL U35 ( .A(n63), .B(n64), .Z(n62) );
  CND2XL U36 ( .A(n55), .B(n53), .Z(n56) );
  CENX1 U37 ( .A(n19), .B(n12), .Z(SUM[25]) );
  CND2XL U38 ( .A(n29), .B(n23), .Z(n19) );
  CND2XL U39 ( .A(n44), .B(n45), .Z(n43) );
  CANR1X1 U40 ( .A(n141), .B(n142), .C(n143), .Z(n136) );
  CND2IXL U41 ( .B(n73), .A(n72), .Z(n74) );
  CND2XL U42 ( .A(n47), .B(n49), .Z(n50) );
  CEOXL U43 ( .A(n107), .B(n108), .Z(SUM[18]) );
  CENX1 U44 ( .A(n20), .B(n5), .Z(SUM[17]) );
  CND2XL U45 ( .A(n91), .B(n14), .Z(n20) );
  CENX1 U46 ( .A(n21), .B(n6), .Z(SUM[13]) );
  CND2XL U47 ( .A(n122), .B(n2), .Z(n21) );
  COND1X1 U48 ( .A(n51), .B(n52), .C(n53), .Z(n46) );
  CIVXL U49 ( .A(n54), .Z(n52) );
  CND2XL U50 ( .A(B[6]), .B(A[6]), .Z(n49) );
  CNR3X1 U51 ( .A(n144), .B(n145), .C(n146), .Z(n143) );
  CNR2XL U52 ( .A(A[6]), .B(B[6]), .Z(n157) );
  CNR2XL U53 ( .A(A[5]), .B(B[5]), .Z(n158) );
  CND2XL U54 ( .A(B[3]), .B(A[3]), .Z(n64) );
  COR2XL U55 ( .A(B[1]), .B(A[1]), .Z(n82) );
  CND2XL U56 ( .A(n71), .B(n72), .Z(n69) );
  CEOXL U57 ( .A(n69), .B(n70), .Z(SUM[31]) );
  CND2XL U58 ( .A(B[0]), .B(A[0]), .Z(n148) );
  CNR2XL U59 ( .A(A[1]), .B(B[1]), .Z(n147) );
  CND2XL U60 ( .A(B[4]), .B(A[4]), .Z(n155) );
  COR2XL U61 ( .A(B[2]), .B(A[2]), .Z(n66) );
  CANR1XL U62 ( .A(n33), .B(n34), .C(n35), .Z(n32) );
  CENX1 U63 ( .A(n32), .B(n31), .Z(SUM[9]) );
  CNR2X1 U64 ( .A(n114), .B(n115), .Z(n120) );
  CENX1 U65 ( .A(n36), .B(n37), .Z(SUM[8]) );
  CANR1XL U66 ( .A(n38), .B(n39), .C(n40), .Z(n36) );
  CND2IX1 U67 ( .B(n85), .A(n72), .Z(n86) );
  CND2XL U68 ( .A(n60), .B(n38), .Z(n34) );
  CNR2X1 U69 ( .A(n114), .B(n115), .Z(n113) );
  CND2X1 U70 ( .A(n125), .B(n126), .Z(n123) );
  CANR1XL U71 ( .A(n118), .B(n33), .C(n115), .Z(n125) );
  CAN4X1 U72 ( .A(n29), .B(n25), .C(n12), .D(n4), .Z(n22) );
  CND3X1 U73 ( .A(n119), .B(n120), .C(n60), .Z(n109) );
  CNR2X1 U74 ( .A(n116), .B(n117), .Z(n111) );
  CND4X1 U75 ( .A(n127), .B(n128), .C(n8), .D(n3), .Z(n115) );
  CND4X1 U76 ( .A(n47), .B(n45), .C(n55), .D(n59), .Z(n118) );
  CNR2IX1 U77 ( .B(n64), .A(n138), .Z(n137) );
  CENX1 U78 ( .A(n56), .B(n54), .Z(SUM[5]) );
  CENX1 U79 ( .A(n9), .B(n1), .Z(SUM[14]) );
  CEOX1 U80 ( .A(n61), .B(n62), .Z(SUM[3]) );
  CANR1XL U81 ( .A(n65), .B(n66), .C(n67), .Z(n61) );
  CND2X1 U82 ( .A(n112), .B(n45), .Z(n33) );
  CND3XL U83 ( .A(n13), .B(n1), .C(n2), .Z(n114) );
  CAN2X1 U84 ( .A(n27), .B(n101), .Z(n25) );
  CENX1 U85 ( .A(n89), .B(n88), .Z(SUM[27]) );
  CEOX1 U86 ( .A(n42), .B(n43), .Z(SUM[7]) );
  CANR1XL U87 ( .A(n46), .B(n47), .C(n48), .Z(n42) );
  CENX1 U88 ( .A(n50), .B(n46), .Z(SUM[6]) );
  CENX1 U89 ( .A(n131), .B(n128), .Z(SUM[10]) );
  CND2XL U90 ( .A(n28), .B(n91), .Z(n107) );
  CEOXL U91 ( .A(n14), .B(n91), .Z(SUM[16]) );
  CENX1 U92 ( .A(n2), .B(n123), .Z(SUM[12]) );
  CEOX1 U93 ( .A(n104), .B(n105), .Z(SUM[19]) );
  CND2XL U94 ( .A(n27), .B(n91), .Z(n104) );
  CENX1 U95 ( .A(n102), .B(n81), .Z(SUM[1]) );
  CND2X1 U96 ( .A(n82), .B(n80), .Z(n102) );
  CENX1 U97 ( .A(n77), .B(n65), .Z(SUM[2]) );
  CND2X1 U98 ( .A(n66), .B(n68), .Z(n77) );
  CNR2IX1 U99 ( .B(n6), .A(n118), .Z(n119) );
  CENX1 U100 ( .A(n93), .B(n92), .Z(SUM[24]) );
  CEOX1 U101 ( .A(n96), .B(n97), .Z(SUM[23]) );
  CND2XL U102 ( .A(n30), .B(n23), .Z(n96) );
  CND2XL U103 ( .A(n76), .B(n72), .Z(n83) );
  CND2X1 U104 ( .A(n10), .B(n72), .Z(n89) );
  CND2X1 U105 ( .A(n10), .B(n88), .Z(n85) );
  CAN2X1 U106 ( .A(n30), .B(n95), .Z(n26) );
  CAN2X1 U107 ( .A(n28), .B(n11), .Z(n27) );
  CAN2X1 U108 ( .A(n14), .B(n5), .Z(n28) );
  CEOXL U109 ( .A(n10), .B(n72), .Z(SUM[26]) );
  CENX1 U110 ( .A(n100), .B(n7), .Z(SUM[21]) );
  CAN2X1 U111 ( .A(n26), .B(n92), .Z(n29) );
  COND2X1 U112 ( .A(n134), .B(n135), .C(n34), .D(n135), .Z(n133) );
  CND2XL U113 ( .A(n3), .B(n8), .Z(n135) );
  COND1XL U114 ( .A(n78), .B(n79), .C(n80), .Z(n65) );
  CND2X1 U115 ( .A(B[1]), .B(A[1]), .Z(n144) );
  CNR2X1 U116 ( .A(A[3]), .B(B[3]), .Z(n145) );
  CNR2IX1 U117 ( .B(B[28]), .A(n85), .Z(n76) );
  COR2X1 U118 ( .A(B[7]), .B(A[7]), .Z(n45) );
  CEOX1 U119 ( .A(n74), .B(n75), .Z(SUM[30]) );
  CEOX1 U120 ( .A(n83), .B(n84), .Z(SUM[29]) );
  CEOX1 U121 ( .A(n86), .B(n87), .Z(SUM[28]) );
  COR2X1 U122 ( .A(B[4]), .B(A[4]), .Z(n59) );
  COR2X1 U123 ( .A(B[5]), .B(A[5]), .Z(n55) );
  CND3X1 U124 ( .A(n152), .B(n153), .C(n154), .Z(n112) );
  CNR2IX1 U125 ( .B(B[30]), .A(n73), .Z(n71) );
  CNR2X1 U126 ( .A(n149), .B(n150), .Z(n141) );
  CNR2XL U127 ( .A(A[3]), .B(B[3]), .Z(n149) );
  CNR2XL U128 ( .A(A[2]), .B(B[2]), .Z(n150) );
  CNR2X1 U129 ( .A(n147), .B(n148), .Z(n142) );
  CND2XL U130 ( .A(B[4]), .B(A[4]), .Z(n58) );
  CND2XL U131 ( .A(B[5]), .B(A[5]), .Z(n53) );
  CND2XL U132 ( .A(B[1]), .B(A[1]), .Z(n80) );
  CND2XL U133 ( .A(B[2]), .B(A[2]), .Z(n68) );
  CAN2X1 U134 ( .A(B[21]), .B(B[22]), .Z(n30) );
  COR2X1 U135 ( .A(B[3]), .B(A[3]), .Z(n63) );
  CNR2X1 U136 ( .A(n157), .B(n158), .Z(n156) );
  CND2X1 U137 ( .A(B[29]), .B(n76), .Z(n73) );
  CND2XL U138 ( .A(B[7]), .B(A[7]), .Z(n44) );
  CND2XL U139 ( .A(B[0]), .B(A[0]), .Z(n103) );
  CND2XL U140 ( .A(A[2]), .B(B[2]), .Z(n140) );
  COR2X1 U141 ( .A(B[6]), .B(A[6]), .Z(n47) );
  CAN2X1 U142 ( .A(n103), .B(n151), .Z(SUM[0]) );
  CND2X1 U143 ( .A(n159), .B(n160), .Z(n151) );
  CIVX2 U144 ( .A(n95), .Z(n97) );
  CIVX2 U145 ( .A(n101), .Z(n105) );
  CIVX2 U146 ( .A(n11), .Z(n108) );
  CIVX2 U147 ( .A(n123), .Z(n122) );
  CIVX2 U148 ( .A(n41), .Z(n39) );
  CIVX2 U149 ( .A(n35), .Z(n37) );
  CIVX2 U150 ( .A(n40), .Z(n134) );
  CND2X2 U151 ( .A(n109), .B(n110), .Z(n91) );
  CIVX2 U152 ( .A(n90), .Z(n88) );
  CIVX2 U153 ( .A(n94), .Z(n92) );
  CIVX2 U154 ( .A(n98), .Z(n95) );
  CIVX2 U155 ( .A(n103), .Z(n81) );
  CIVX2 U156 ( .A(n106), .Z(n101) );
  CIVX2 U157 ( .A(n132), .Z(n127) );
  CIVX2 U158 ( .A(n124), .Z(n128) );
  CIVX2 U159 ( .A(B[28]), .Z(n87) );
  CIVX2 U160 ( .A(B[29]), .Z(n84) );
  CIVX2 U161 ( .A(B[30]), .Z(n75) );
  CIVX2 U162 ( .A(B[31]), .Z(n70) );
  CIVX2 U163 ( .A(n8), .Z(n31) );
  CIVX2 U164 ( .A(n3), .Z(n35) );
  CIVX2 U165 ( .A(n49), .Z(n48) );
  CIVX2 U166 ( .A(n55), .Z(n51) );
  CIVX2 U167 ( .A(n59), .Z(n57) );
  CIVX2 U168 ( .A(n68), .Z(n67) );
  CIVX2 U169 ( .A(n81), .Z(n79) );
  CIVX2 U170 ( .A(n82), .Z(n78) );
  CIVX2 U171 ( .A(B[24]), .Z(n94) );
  CIVX2 U172 ( .A(B[23]), .Z(n98) );
  CIVX2 U173 ( .A(n7), .Z(n99) );
  CIVX2 U174 ( .A(n23), .Z(n100) );
  CIVX2 U175 ( .A(B[19]), .Z(n106) );
  CND3X1 U176 ( .A(n111), .B(n112), .C(n113), .Z(n110) );
  CIVX2 U177 ( .A(n6), .Z(n117) );
  CIVX2 U178 ( .A(n45), .Z(n116) );
  CIVX2 U179 ( .A(n1), .Z(n121) );
  CIVX2 U180 ( .A(n60), .Z(n41) );
  CIVX2 U181 ( .A(n128), .Z(n130) );
  CIVX2 U182 ( .A(B[11]), .Z(n132) );
  CIVX2 U183 ( .A(B[10]), .Z(n124) );
  CIVX2 U184 ( .A(n133), .Z(n131) );
  CIVX2 U185 ( .A(n118), .Z(n38) );
  CND2X2 U186 ( .A(n136), .B(n137), .Z(n60) );
  CIVX2 U187 ( .A(n63), .Z(n139) );
  CIVX2 U188 ( .A(n33), .Z(n40) );
  CND2IX1 U189 ( .B(n155), .A(n156), .Z(n154) );
  COND3X1 U190 ( .A(A[6]), .B(B[6]), .C(A[5]), .D(B[5]), .Z(n153) );
  CAN2X1 U191 ( .A(n44), .B(n49), .Z(n152) );
  CIVX2 U192 ( .A(A[0]), .Z(n160) );
  CIVX2 U193 ( .A(B[0]), .Z(n159) );
endmodule


module nios_2_DW01_cmp6_2 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255;

  CANR11X1 U1 ( .A(n76), .B(n77), .C(n78), .D(n79), .Z(n75) );
  CNR3X2 U2 ( .A(n206), .B(n207), .C(n208), .Z(n193) );
  CIVXL U3 ( .A(n178), .Z(n1) );
  CND2X1 U4 ( .A(n103), .B(n104), .Z(n100) );
  CNR3X1 U5 ( .A(n213), .B(n214), .C(n7), .Z(n212) );
  CIVX2 U6 ( .A(A[14]), .Z(n167) );
  CNR2X2 U7 ( .A(n105), .B(n106), .Z(n98) );
  CIVX1 U8 ( .A(n63), .Z(n106) );
  CNR2IXL U9 ( .B(n160), .A(n191), .Z(n185) );
  CIVXL U10 ( .A(A[29]), .Z(n251) );
  CNR2X1 U11 ( .A(n242), .B(n243), .Z(n237) );
  CND2IXL U12 ( .B(A[30]), .A(B[30]), .Z(n250) );
  CNR3X2 U13 ( .A(n100), .B(n66), .C(n67), .Z(n99) );
  CND2X1 U14 ( .A(A[11]), .B(n101), .Z(n42) );
  CIVX1 U15 ( .A(n95), .Z(n93) );
  CIVX1 U16 ( .A(n42), .Z(n67) );
  CNR2XL U17 ( .A(B[14]), .B(n203), .Z(n202) );
  CIVX1 U18 ( .A(A[4]), .Z(n188) );
  CND3XL U19 ( .A(n181), .B(n182), .C(n183), .Z(n175) );
  CND2XL U20 ( .A(B[8]), .B(n157), .Z(n56) );
  CIVXL U21 ( .A(n167), .Z(n2) );
  CND2X1 U22 ( .A(B[10]), .B(n156), .Z(n72) );
  CIVX1 U23 ( .A(n43), .Z(n66) );
  CIVX2 U24 ( .A(A[24]), .Z(n171) );
  CND2X1 U25 ( .A(A[24]), .B(n230), .Z(n124) );
  CIVXL U26 ( .A(n248), .Z(n13) );
  CND4XL U27 ( .A(n113), .B(n250), .C(n249), .D(n122), .Z(n248) );
  CNR2IX2 U28 ( .B(n15), .A(n12), .Z(GT) );
  CENX1 U29 ( .A(B[31]), .B(A[31]), .Z(n112) );
  CND4X1 U30 ( .A(A[26]), .B(n129), .C(n122), .D(n252), .Z(n134) );
  CND2X2 U31 ( .A(B[27]), .B(n253), .Z(n129) );
  CIVXL U32 ( .A(B[24]), .Z(n230) );
  CIVXL U33 ( .A(B[1]), .Z(n178) );
  CIVXL U34 ( .A(n21), .Z(n137) );
  CND3X1 U35 ( .A(n126), .B(n130), .C(n121), .Z(n169) );
  CND4XL U36 ( .A(n26), .B(n10), .C(n27), .D(n28), .Z(n24) );
  CNR2XL U37 ( .A(B[18]), .B(n209), .Z(n208) );
  CIVX1 U38 ( .A(A[23]), .Z(n172) );
  CND4XL U39 ( .A(n45), .B(n2), .C(n82), .D(n202), .Z(n194) );
  CIVXL U40 ( .A(A[1]), .Z(n189) );
  CNR2XL U41 ( .A(A[1]), .B(n178), .Z(n191) );
  COND2XL U42 ( .A(A[1]), .B(n178), .C(A[0]), .D(n179), .Z(n177) );
  CIVXL U43 ( .A(A[19]), .Z(n174) );
  CND2X2 U44 ( .A(A[19]), .B(n210), .Z(n53) );
  CND2IXL U45 ( .B(A[20]), .A(B[20]), .Z(n173) );
  CND2IXL U46 ( .B(A[20]), .A(B[20]), .Z(n46) );
  CIVXL U47 ( .A(A[7]), .Z(n158) );
  CND2X2 U48 ( .A(A[7]), .B(n244), .Z(n103) );
  CNR2XL U49 ( .A(n58), .B(n59), .Z(n32) );
  CND3X2 U50 ( .A(n140), .B(n141), .C(n142), .Z(n86) );
  CIVX1 U51 ( .A(A[21]), .Z(n219) );
  CIVXL U52 ( .A(A[18]), .Z(n52) );
  CIVXL U53 ( .A(A[18]), .Z(n209) );
  CIVXL U54 ( .A(A[6]), .Z(n161) );
  CND2X1 U55 ( .A(A[6]), .B(n241), .Z(n104) );
  CND2IXL U56 ( .B(B[12]), .A(A[12]), .Z(n44) );
  CND2IXL U57 ( .B(B[13]), .A(A[13]), .Z(n236) );
  CND2IXL U58 ( .B(A[13]), .A(B[13]), .Z(n81) );
  CIVXL U59 ( .A(A[13]), .Z(n71) );
  CIVXL U60 ( .A(A[11]), .Z(n247) );
  CND2X1 U61 ( .A(n65), .B(n99), .Z(n3) );
  CND2X2 U62 ( .A(n98), .B(n4), .Z(n97) );
  CIVX1 U63 ( .A(n3), .Z(n4) );
  CND3X1 U64 ( .A(n41), .B(n72), .C(n8), .Z(n65) );
  CIVX1 U65 ( .A(A[9]), .Z(n166) );
  CND2X2 U66 ( .A(B[17]), .B(n205), .Z(n82) );
  CND3XL U67 ( .A(B[18]), .B(n52), .C(n53), .Z(n28) );
  CIVXL U68 ( .A(B[15]), .Z(n200) );
  CND2IXL U69 ( .B(A[18]), .A(B[18]), .Z(n165) );
  CNR3X1 U70 ( .A(n47), .B(n30), .C(n215), .Z(n213) );
  CNR2X1 U71 ( .A(n22), .B(n233), .Z(n136) );
  CND2X1 U72 ( .A(n11), .B(n12), .Z(NE) );
  CND2X2 U73 ( .A(B[28]), .B(n255), .Z(n122) );
  CND4XL U74 ( .A(n91), .B(n96), .C(n159), .D(n160), .Z(n154) );
  CNR2X1 U75 ( .A(n163), .B(n164), .Z(n152) );
  CNR2X1 U76 ( .A(n14), .B(n86), .Z(n139) );
  CNR2X1 U77 ( .A(n29), .B(n30), .Z(n27) );
  CNR2X1 U78 ( .A(n215), .B(n216), .Z(n214) );
  CNR2X1 U79 ( .A(n35), .B(n36), .Z(n34) );
  CND2XL U80 ( .A(n39), .B(n40), .Z(n38) );
  CNR2IXL U81 ( .B(n60), .A(n57), .Z(n59) );
  CNR2XL U82 ( .A(n72), .B(n57), .Z(n58) );
  CAN3XL U83 ( .A(n93), .B(n44), .C(n40), .Z(n6) );
  CNR2IX1 U84 ( .B(A[9]), .A(B[9]), .Z(n9) );
  CND4X1 U85 ( .A(n80), .B(n95), .C(n54), .D(n41), .Z(n163) );
  CNR2XL U86 ( .A(B[12]), .B(n70), .Z(n69) );
  COND2XL U87 ( .A(n1), .B(n189), .C(B[0]), .D(n190), .Z(n186) );
  CND2X1 U88 ( .A(B[19]), .B(n174), .Z(n31) );
  CND4XL U89 ( .A(n80), .B(n81), .C(n82), .D(n83), .Z(n79) );
  CNR2XL U90 ( .A(n25), .B(n184), .Z(n138) );
  CND2XL U91 ( .A(n84), .B(n85), .Z(n184) );
  CNR2IXL U92 ( .B(n111), .A(n7), .Z(n110) );
  CND3XL U93 ( .A(n61), .B(n56), .C(n72), .Z(n155) );
  CND2XL U94 ( .A(n90), .B(n31), .Z(n89) );
  CAN3XL U95 ( .A(n134), .B(n133), .C(n5), .Z(n107) );
  CAN2XL U96 ( .A(n131), .B(n132), .Z(n5) );
  CNR2XL U97 ( .A(n145), .B(n146), .Z(n187) );
  CND2X1 U98 ( .A(B[22]), .B(n218), .Z(n26) );
  CNR2IXL U99 ( .B(A[31]), .A(B[31]), .Z(n7) );
  CNR2IX1 U100 ( .B(A[2]), .A(n146), .Z(n143) );
  CND2XL U101 ( .A(A[13]), .B(n94), .Z(n40) );
  CND2X1 U102 ( .A(B[29]), .B(n251), .Z(n113) );
  CND4XL U103 ( .A(n90), .B(n31), .C(n173), .D(n82), .Z(n168) );
  CNR2XL U104 ( .A(B[17]), .B(n205), .Z(n207) );
  CNR2XL U105 ( .A(B[3]), .B(n149), .Z(n147) );
  CND2IXL U106 ( .B(A[16]), .A(B[16]), .Z(n183) );
  CENXL U107 ( .A(B[31]), .B(A[31]), .Z(n249) );
  CND2X1 U108 ( .A(A[21]), .B(n217), .Z(n216) );
  COND1X1 U109 ( .A(n17), .B(n18), .C(n19), .Z(n16) );
  CND2IXL U110 ( .B(B[4]), .A(A[4]), .Z(n84) );
  CND2IXL U111 ( .B(A[4]), .A(B[4]), .Z(n182) );
  CNR2X1 U112 ( .A(n20), .B(n21), .Z(n19) );
  CND3XL U113 ( .A(n32), .B(n33), .C(n34), .Z(n18) );
  CANR3X1 U114 ( .A(n48), .B(n49), .C(n50), .D(n51), .Z(n33) );
  CNR2X1 U115 ( .A(n54), .B(n55), .Z(n50) );
  CND4X1 U116 ( .A(n150), .B(n151), .C(n152), .D(n153), .Z(n14) );
  CNR2X1 U117 ( .A(n168), .B(n169), .Z(n151) );
  CNR3X1 U118 ( .A(n175), .B(n176), .C(n177), .Z(n150) );
  CNR2X1 U119 ( .A(n154), .B(n155), .Z(n153) );
  CANR1X1 U120 ( .A(n87), .B(n88), .C(n89), .Z(n74) );
  CANR1X1 U121 ( .A(n88), .B(n92), .C(n6), .Z(n73) );
  CND2X1 U122 ( .A(n147), .B(n148), .Z(n140) );
  CNR2X1 U123 ( .A(n8), .B(n9), .Z(n141) );
  CND2X1 U124 ( .A(n143), .B(n144), .Z(n142) );
  CND2XL U125 ( .A(n13), .B(n76), .Z(n233) );
  CAN2X1 U126 ( .A(n84), .B(n85), .Z(n78) );
  CND3XL U127 ( .A(n114), .B(n115), .C(n116), .Z(n108) );
  CND3XL U128 ( .A(n123), .B(n124), .C(n125), .Z(n115) );
  CANR1XL U129 ( .A(n123), .B(n127), .C(n128), .Z(n114) );
  CNR3XL U130 ( .A(n117), .B(n118), .C(n119), .Z(n116) );
  CND3XL U131 ( .A(n42), .B(n43), .C(n44), .Z(n37) );
  CNR2IXL U132 ( .B(n13), .A(n14), .Z(n11) );
  CND2X1 U133 ( .A(n211), .B(n212), .Z(n21) );
  CNR2X1 U134 ( .A(n220), .B(n221), .Z(n211) );
  CNR2X1 U135 ( .A(n37), .B(n38), .Z(n36) );
  CND3XL U136 ( .A(n45), .B(n26), .C(n10), .Z(n35) );
  CND2X1 U137 ( .A(n9), .B(n72), .Z(n63) );
  CND2X1 U138 ( .A(n133), .B(n134), .Z(n22) );
  CND2X1 U139 ( .A(n111), .B(n131), .Z(n221) );
  CND2X1 U140 ( .A(n129), .B(n120), .Z(n176) );
  CENX1 U141 ( .A(B[16]), .B(A[16]), .Z(n45) );
  COND2XL U142 ( .A(B[13]), .B(n71), .C(B[12]), .D(n70), .Z(n105) );
  CND4X1 U143 ( .A(n62), .B(n63), .C(n64), .D(n65), .Z(n57) );
  CNR2X1 U144 ( .A(n68), .B(n69), .Z(n62) );
  CNR2X1 U145 ( .A(n66), .B(n67), .Z(n64) );
  CNR2XL U146 ( .A(B[13]), .B(n71), .Z(n68) );
  CNR2X1 U147 ( .A(n231), .B(n232), .Z(n224) );
  CNR2X1 U148 ( .A(n226), .B(n227), .Z(n225) );
  CNR2X1 U149 ( .A(B[23]), .B(n172), .Z(n232) );
  CND4X1 U150 ( .A(n193), .B(n194), .C(n195), .D(n196), .Z(n25) );
  CND2XL U151 ( .A(n197), .B(n82), .Z(n196) );
  CND3X1 U152 ( .A(A[30]), .B(n223), .C(n112), .Z(n111) );
  CND3X1 U153 ( .A(n185), .B(n186), .C(n187), .Z(n85) );
  CNR2X1 U154 ( .A(n239), .B(n240), .Z(n238) );
  CNR2XL U155 ( .A(B[5]), .B(n162), .Z(n239) );
  CNR2XL U156 ( .A(B[12]), .B(n70), .Z(n246) );
  CNR2X1 U157 ( .A(B[2]), .B(n145), .Z(n144) );
  CND2X1 U158 ( .A(B[9]), .B(n166), .Z(n41) );
  CND3XL U159 ( .A(n83), .B(n165), .C(n81), .Z(n164) );
  CNR2XL U160 ( .A(B[10]), .B(n156), .Z(n243) );
  CNR2XL U161 ( .A(B[11]), .B(n247), .Z(n245) );
  CNR2XL U162 ( .A(B[16]), .B(n198), .Z(n197) );
  CND2X1 U163 ( .A(B[21]), .B(n219), .Z(n90) );
  CND2X1 U164 ( .A(B[15]), .B(n204), .Z(n83) );
  CNR2IX1 U165 ( .B(A[8]), .A(B[8]), .Z(n8) );
  CND2X1 U166 ( .A(A[29]), .B(n222), .Z(n131) );
  CND4X1 U167 ( .A(n235), .B(n236), .C(n237), .D(n238), .Z(n234) );
  CNR2X1 U168 ( .A(n245), .B(n246), .Z(n235) );
  CND2X1 U169 ( .A(B[26]), .B(n170), .Z(n121) );
  CND2X1 U170 ( .A(B[2]), .B(n192), .Z(n160) );
  CND2X1 U171 ( .A(A[28]), .B(n228), .Z(n132) );
  CND2X1 U172 ( .A(B[25]), .B(n180), .Z(n120) );
  CND2X1 U173 ( .A(B[4]), .B(n188), .Z(n148) );
  CND2X1 U174 ( .A(B[3]), .B(n149), .Z(n159) );
  CND2X1 U175 ( .A(A[10]), .B(n102), .Z(n43) );
  CND2X1 U176 ( .A(B[24]), .B(n171), .Z(n130) );
  CND2X1 U177 ( .A(n254), .B(n122), .Z(n133) );
  CNR2XL U178 ( .A(B[27]), .B(n253), .Z(n254) );
  CND2X1 U179 ( .A(B[14]), .B(n167), .Z(n80) );
  CND3XL U180 ( .A(n112), .B(n250), .C(n113), .Z(n109) );
  CND2X1 U181 ( .A(B[7]), .B(n158), .Z(n61) );
  CND2X1 U182 ( .A(B[23]), .B(n172), .Z(n126) );
  CND2X1 U183 ( .A(B[5]), .B(n162), .Z(n91) );
  CND4X1 U184 ( .A(n136), .B(n137), .C(n138), .D(n139), .Z(n135) );
  CND2X1 U185 ( .A(A[25]), .B(n229), .Z(n123) );
  CAN2X1 U186 ( .A(n46), .B(n47), .Z(n10) );
  CND3XL U187 ( .A(n45), .B(A[15]), .C(n199), .Z(n195) );
  CNR2IX1 U188 ( .B(n200), .A(n201), .Z(n199) );
  CIVX1 U189 ( .A(B[28]), .Z(n228) );
  CND2X1 U190 ( .A(B[6]), .B(n161), .Z(n96) );
  CNR2XL U191 ( .A(B[22]), .B(n218), .Z(n231) );
  CND2IXL U192 ( .B(A[22]), .A(B[22]), .Z(n181) );
  CIVX2 U193 ( .A(n16), .Z(n12) );
  CND2IX1 U194 ( .B(n22), .A(n23), .Z(n20) );
  CND2IX1 U195 ( .B(n24), .A(n25), .Z(n23) );
  CIVX2 U196 ( .A(n31), .Z(n29) );
  CIVX2 U197 ( .A(n41), .Z(n39) );
  CIVX2 U198 ( .A(n28), .Z(n51) );
  CIVX2 U199 ( .A(n40), .Z(n55) );
  CIVX2 U200 ( .A(n56), .Z(n49) );
  CIVX2 U201 ( .A(n57), .Z(n48) );
  CIVX2 U202 ( .A(n61), .Z(n60) );
  CND3X1 U203 ( .A(n75), .B(n74), .C(n73), .Z(n17) );
  CIVX2 U204 ( .A(n86), .Z(n77) );
  CIVX2 U205 ( .A(n91), .Z(n87) );
  CIVX2 U206 ( .A(B[13]), .Z(n94) );
  CIVX2 U207 ( .A(n96), .Z(n92) );
  CIVX2 U208 ( .A(n97), .Z(n88) );
  CIVX2 U209 ( .A(B[11]), .Z(n101) );
  CIVX2 U210 ( .A(B[10]), .Z(n102) );
  COND4CX1 U211 ( .A(n107), .B(n108), .C(n109), .D(n110), .Z(n15) );
  CIVX2 U212 ( .A(n120), .Z(n119) );
  CIVX2 U213 ( .A(n121), .Z(n118) );
  CIVX2 U214 ( .A(n122), .Z(n117) );
  CIVX2 U215 ( .A(n126), .Z(n125) );
  CIVX2 U216 ( .A(n129), .Z(n128) );
  CIVX2 U217 ( .A(n130), .Z(n127) );
  CIVX2 U218 ( .A(n135), .Z(EQ) );
  CIVX2 U219 ( .A(A[8]), .Z(n157) );
  CND2IX1 U220 ( .B(A[12]), .A(B[12]), .Z(n54) );
  CND2IX1 U221 ( .B(A[11]), .A(B[11]), .Z(n95) );
  CIVX2 U222 ( .A(A[26]), .Z(n170) );
  CIVX2 U223 ( .A(B[0]), .Z(n179) );
  CIVX2 U224 ( .A(A[25]), .Z(n180) );
  CIVX2 U225 ( .A(n159), .Z(n146) );
  CIVX2 U226 ( .A(A[3]), .Z(n149) );
  CIVX2 U227 ( .A(n148), .Z(n145) );
  CIVX2 U228 ( .A(A[0]), .Z(n190) );
  CIVX2 U229 ( .A(A[2]), .Z(n192) );
  CIVX2 U230 ( .A(A[16]), .Z(n198) );
  CIVX2 U231 ( .A(n82), .Z(n201) );
  CIVX2 U232 ( .A(n83), .Z(n203) );
  CIVX2 U233 ( .A(A[15]), .Z(n204) );
  CIVX2 U234 ( .A(A[17]), .Z(n205) );
  CIVX2 U235 ( .A(n53), .Z(n206) );
  CIVX2 U236 ( .A(B[19]), .Z(n210) );
  CIVX2 U237 ( .A(B[21]), .Z(n217) );
  CIVX2 U238 ( .A(n26), .Z(n215) );
  CIVX2 U239 ( .A(n90), .Z(n30) );
  CND2IX1 U240 ( .B(B[20]), .A(A[20]), .Z(n47) );
  CIVX2 U241 ( .A(B[29]), .Z(n222) );
  CIVX2 U242 ( .A(B[30]), .Z(n223) );
  CND3X1 U243 ( .A(n224), .B(n124), .C(n225), .Z(n220) );
  CIVX2 U244 ( .A(n132), .Z(n227) );
  CIVX2 U245 ( .A(n123), .Z(n226) );
  CIVX2 U246 ( .A(B[25]), .Z(n229) );
  CIVX2 U247 ( .A(A[22]), .Z(n218) );
  CIVX2 U248 ( .A(n234), .Z(n76) );
  CIVX2 U249 ( .A(n104), .Z(n240) );
  CIVX2 U250 ( .A(B[6]), .Z(n241) );
  CIVX2 U251 ( .A(A[5]), .Z(n162) );
  CIVX2 U252 ( .A(A[10]), .Z(n156) );
  CIVX2 U253 ( .A(n103), .Z(n242) );
  CIVX2 U254 ( .A(B[7]), .Z(n244) );
  CIVX2 U255 ( .A(A[12]), .Z(n70) );
  CIVX2 U256 ( .A(B[26]), .Z(n252) );
  CIVX2 U257 ( .A(A[28]), .Z(n255) );
  CIVX2 U258 ( .A(A[27]), .Z(n253) );
endmodule


module nios_2_DW01_sub_3 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357;

  CND2X1 U3 ( .A(A[20]), .B(n206), .Z(n187) );
  CENX1 U4 ( .A(n133), .B(n9), .Z(DIFF[28]) );
  CAN3X1 U5 ( .A(n96), .B(n95), .C(n12), .Z(n1) );
  CNIVX1 U6 ( .A(n93), .Z(n2) );
  CIVXL U7 ( .A(B[8]), .Z(n330) );
  CIVX1 U8 ( .A(n110), .Z(n18) );
  CIVXL U9 ( .A(n189), .Z(n3) );
  CIVX2 U10 ( .A(n3), .Z(n4) );
  CND2IX2 U11 ( .B(A[21]), .A(B[21]), .Z(n196) );
  CIVX2 U12 ( .A(n194), .Z(n189) );
  CND2IX2 U13 ( .B(A[20]), .A(B[20]), .Z(n195) );
  CNIVX1 U14 ( .A(n116), .Z(n5) );
  CIVX2 U15 ( .A(n137), .Z(n116) );
  CIVXL U16 ( .A(n187), .Z(n198) );
  CIVX1 U17 ( .A(n273), .Z(n302) );
  CIVXL U18 ( .A(B[24]), .Z(n175) );
  CND2X1 U19 ( .A(B[24]), .B(n176), .Z(n147) );
  CND3X1 U20 ( .A(n143), .B(n144), .C(n145), .Z(n132) );
  CIVX2 U21 ( .A(n317), .Z(n6) );
  CND2XL U22 ( .A(n167), .B(n168), .Z(n183) );
  CNIVXL U23 ( .A(n60), .Z(n7) );
  CENXL U24 ( .A(n286), .B(n287), .Z(DIFF[15]) );
  CND2XL U25 ( .A(n130), .B(n126), .Z(n136) );
  CAN2X2 U26 ( .A(n113), .B(n114), .Z(n39) );
  CIVX1 U27 ( .A(n261), .Z(n334) );
  CIVX1 U28 ( .A(n49), .Z(n328) );
  CENXL U29 ( .A(n190), .B(n191), .Z(DIFF[22]) );
  CIVXL U30 ( .A(n245), .Z(n8) );
  CND2IX2 U31 ( .B(n30), .A(n315), .Z(n245) );
  CENXL U32 ( .A(B[28]), .B(A[28]), .Z(n9) );
  CIVX2 U33 ( .A(n170), .Z(n10) );
  CIVXL U34 ( .A(n170), .Z(n119) );
  CND2IX1 U35 ( .B(n303), .A(n304), .Z(n273) );
  CENXL U36 ( .A(n139), .B(n43), .Z(DIFF[27]) );
  CDLY1XL U37 ( .A(n312), .Z(n15) );
  CND2XL U38 ( .A(n94), .B(n92), .Z(n11) );
  CIVX2 U39 ( .A(n11), .Z(n12) );
  CND2X2 U40 ( .A(n101), .B(n88), .Z(n94) );
  CNR2IX2 U41 ( .B(n118), .A(n164), .Z(n163) );
  CND3X1 U42 ( .A(n273), .B(n274), .C(n270), .Z(n237) );
  CND2X1 U43 ( .A(A[27]), .B(n141), .Z(n129) );
  CND2X1 U44 ( .A(A[18]), .B(n225), .Z(n210) );
  CIVX2 U45 ( .A(n305), .Z(n318) );
  CIVX2 U46 ( .A(n245), .Z(n260) );
  CND4X1 U47 ( .A(n340), .B(n215), .C(n80), .D(n82), .Z(n249) );
  CND2X1 U48 ( .A(B[9]), .B(n329), .Z(n50) );
  CNR2IXL U49 ( .B(n130), .A(n131), .Z(n142) );
  CNR2IXL U50 ( .B(n221), .A(n227), .Z(n226) );
  COND1X1 U51 ( .A(n253), .B(n288), .C(n283), .Z(n287) );
  CND2XL U52 ( .A(n313), .B(n319), .Z(n322) );
  CAN2X1 U53 ( .A(n230), .B(n231), .Z(n13) );
  CIVXL U54 ( .A(A[5]), .Z(n336) );
  CIVX1 U55 ( .A(B[3]), .Z(n339) );
  CND2XL U56 ( .A(B[4]), .B(n335), .Z(n73) );
  CANR1X1 U57 ( .A(n59), .B(n7), .C(n61), .Z(n56) );
  CND2X2 U58 ( .A(B[6]), .B(n352), .Z(n60) );
  CIVXL U59 ( .A(n332), .Z(n14) );
  CIVX3 U60 ( .A(n268), .Z(n250) );
  CIVX1 U61 ( .A(n26), .Z(n204) );
  COND1X1 U62 ( .A(n316), .B(n52), .C(n55), .Z(n49) );
  CND2X2 U63 ( .A(n24), .B(n2), .Z(n35) );
  CND2X1 U64 ( .A(B[2]), .B(n341), .Z(n80) );
  CND3X2 U65 ( .A(n220), .B(n221), .C(n222), .Z(n209) );
  CENXL U66 ( .A(n177), .B(n178), .Z(DIFF[23]) );
  CIVX1 U67 ( .A(n58), .Z(n333) );
  CND2X1 U68 ( .A(n55), .B(n51), .Z(n306) );
  CND2XL U69 ( .A(A[13]), .B(n299), .Z(n16) );
  CND2IX1 U70 ( .B(n17), .A(n281), .Z(n275) );
  CNR3X1 U71 ( .A(n250), .B(n280), .C(n253), .Z(n17) );
  CND2XL U72 ( .A(n299), .B(A[13]), .Z(n280) );
  CND2IX2 U73 ( .B(A[15]), .A(B[15]), .Z(n268) );
  CNR2IXL U74 ( .B(n81), .A(n251), .Z(n248) );
  CENXL U75 ( .A(n201), .B(n202), .Z(DIFF[21]) );
  CIVX2 U76 ( .A(n110), .Z(n161) );
  CIVX1 U77 ( .A(B[13]), .Z(n299) );
  CIVX2 U78 ( .A(n325), .Z(n324) );
  CENXL U79 ( .A(n90), .B(n19), .Z(DIFF[29]) );
  CEOXL U80 ( .A(B[29]), .B(A[29]), .Z(n19) );
  COND4CXL U81 ( .A(n160), .B(n161), .C(n162), .D(n163), .Z(n20) );
  COND4CXL U82 ( .A(n160), .B(n161), .C(n162), .D(n163), .Z(n23) );
  CND2X2 U83 ( .A(n90), .B(n47), .Z(n87) );
  CND3X2 U84 ( .A(n38), .B(n100), .C(n103), .Z(n90) );
  COND1XL U85 ( .A(n14), .B(n316), .C(n55), .Z(n21) );
  COND4CX1 U86 ( .A(n160), .B(n18), .C(n162), .D(n163), .Z(n22) );
  COND4CX1 U87 ( .A(n160), .B(n161), .C(n162), .D(n163), .Z(n134) );
  CND2IX2 U88 ( .B(n2), .A(n1), .Z(n36) );
  CAOR1X1 U89 ( .A(n147), .B(n22), .C(n153), .Z(n44) );
  CND4X1 U90 ( .A(n96), .B(n94), .C(n92), .D(n95), .Z(n24) );
  CIVX1 U91 ( .A(n277), .Z(n276) );
  CANR1XL U92 ( .A(n248), .B(n249), .C(n250), .Z(n241) );
  CND2IXL U93 ( .B(B[11]), .A(A[11]), .Z(n313) );
  CIVXL U94 ( .A(B[11]), .Z(n314) );
  CENXL U95 ( .A(n25), .B(n41), .Z(DIFF[18]) );
  CAN2XL U96 ( .A(n210), .B(n222), .Z(n25) );
  COR2XL U97 ( .A(n355), .B(B[10]), .Z(n312) );
  COND1X1 U98 ( .A(n173), .B(n161), .C(n160), .Z(n26) );
  COND1X1 U99 ( .A(n173), .B(n18), .C(n160), .Z(n182) );
  CIVXL U100 ( .A(n205), .Z(n27) );
  CIVX2 U101 ( .A(B[21]), .Z(n205) );
  CIVX2 U102 ( .A(n98), .Z(n97) );
  CIVX1 U103 ( .A(B[7]), .Z(n347) );
  CND2X1 U104 ( .A(A[14]), .B(n294), .Z(n283) );
  CIVXL U105 ( .A(A[14]), .Z(n295) );
  CND2X1 U106 ( .A(n310), .B(A[9]), .Z(n51) );
  CENXL U107 ( .A(n291), .B(n289), .Z(DIFF[14]) );
  CIVX1 U108 ( .A(n289), .Z(n288) );
  COND1X2 U109 ( .A(n34), .B(n52), .C(n302), .Z(n298) );
  CNR2X2 U110 ( .A(n275), .B(n276), .Z(n236) );
  CIVXL U111 ( .A(B[16]), .Z(n284) );
  CND2X1 U112 ( .A(A[15]), .B(n290), .Z(n244) );
  CND2X1 U113 ( .A(A[8]), .B(n330), .Z(n55) );
  CIVXL U114 ( .A(n37), .Z(n28) );
  CIVXL U115 ( .A(n28), .Z(n29) );
  CIVXL U116 ( .A(B[15]), .Z(n290) );
  CND2XL U117 ( .A(n215), .B(n107), .Z(n212) );
  CND2IXL U118 ( .B(B[1]), .A(A[1]), .Z(n107) );
  CND2IXL U119 ( .B(B[1]), .A(A[1]), .Z(n343) );
  CND2X2 U120 ( .A(n126), .B(n138), .Z(n137) );
  CND2X1 U121 ( .A(n54), .B(n50), .Z(n30) );
  CIVXL U122 ( .A(n50), .Z(n317) );
  CNR2XL U123 ( .A(n310), .B(A[9]), .Z(n309) );
  CND2X2 U124 ( .A(B[14]), .B(n295), .Z(n272) );
  CND2IX1 U125 ( .B(B[17]), .A(A[17]), .Z(n228) );
  CIVX1 U126 ( .A(B[2]), .Z(n345) );
  CIVX1 U127 ( .A(n267), .Z(n265) );
  CIVX2 U128 ( .A(n298), .Z(n297) );
  CNR2X1 U129 ( .A(n255), .B(n256), .Z(n31) );
  CANR1X1 U130 ( .A(n138), .B(n23), .C(n142), .Z(n139) );
  CENXL U131 ( .A(n159), .B(n22), .Z(DIFF[24]) );
  CNR2X2 U132 ( .A(n255), .B(n256), .Z(n238) );
  CND2X1 U133 ( .A(n86), .B(n85), .Z(n32) );
  CND2X2 U134 ( .A(n87), .B(n33), .Z(n84) );
  CIVX2 U135 ( .A(n32), .Z(n33) );
  CND2X1 U136 ( .A(n91), .B(n89), .Z(n86) );
  CIVXL U137 ( .A(n8), .Z(n34) );
  CND2X2 U138 ( .A(n116), .B(n117), .Z(n115) );
  CND2X1 U139 ( .A(A[24]), .B(n175), .Z(n158) );
  CIVXL U140 ( .A(A[24]), .Z(n176) );
  CIVXL U141 ( .A(n195), .Z(n203) );
  CND2XL U142 ( .A(n209), .B(n210), .Z(n219) );
  CND3X1 U143 ( .A(n261), .B(n262), .C(n58), .Z(n257) );
  CENX1 U144 ( .A(n150), .B(n151), .Z(DIFF[26]) );
  CND2XL U145 ( .A(n208), .B(n124), .Z(n216) );
  CND2X2 U146 ( .A(B[19]), .B(n218), .Z(n208) );
  COND1X1 U147 ( .A(n234), .B(n161), .C(n229), .Z(n233) );
  CENX1 U148 ( .A(n233), .B(n232), .Z(DIFF[17]) );
  CIVX3 U149 ( .A(n272), .Z(n253) );
  CND2X1 U150 ( .A(n282), .B(n268), .Z(n281) );
  CND2IX1 U151 ( .B(A[17]), .A(B[17]), .Z(n231) );
  CNR2X2 U152 ( .A(n250), .B(n253), .Z(n262) );
  COND1X1 U153 ( .A(n318), .B(n324), .C(n15), .Z(n323) );
  CND2X2 U154 ( .A(n36), .B(n35), .Z(DIFF[30]) );
  CND4X1 U155 ( .A(n31), .B(n236), .C(n237), .D(n239), .Z(n37) );
  CND4X2 U156 ( .A(n236), .B(n238), .C(n237), .D(n239), .Z(n110) );
  CND2IXL U157 ( .B(A[21]), .A(n27), .Z(n197) );
  CANR11X2 U158 ( .A(n242), .B(n240), .C(n241), .D(n243), .Z(n239) );
  CIVX1 U159 ( .A(n244), .Z(n243) );
  CNR3X1 U160 ( .A(n245), .B(n246), .C(n247), .Z(n242) );
  CIVX1 U161 ( .A(B[9]), .Z(n310) );
  COND1X1 U162 ( .A(n64), .B(n65), .C(n66), .Z(n59) );
  CIVX1 U163 ( .A(n69), .Z(n65) );
  CNR2IX4 U164 ( .B(n124), .A(n174), .Z(n160) );
  CIVXL U165 ( .A(B[22]), .Z(n199) );
  CND2XL U166 ( .A(n228), .B(n231), .Z(n232) );
  CND3X1 U167 ( .A(n152), .B(n145), .C(n143), .Z(n151) );
  CND2XL U168 ( .A(n143), .B(n148), .Z(n155) );
  CIVX1 U169 ( .A(B[19]), .Z(n217) );
  COND4CX1 U170 ( .A(n109), .B(n37), .C(n111), .D(n112), .Z(n38) );
  CND3X1 U171 ( .A(n120), .B(n121), .C(n114), .Z(n111) );
  CNR2X2 U172 ( .A(n39), .B(n115), .Z(n112) );
  CNR2IX2 U173 ( .B(n118), .A(n10), .Z(n113) );
  CND2X2 U174 ( .A(n165), .B(n166), .Z(n114) );
  COND4CX1 U175 ( .A(n109), .B(n37), .C(n111), .D(n112), .Z(n98) );
  CEOX1 U176 ( .A(n204), .B(n40), .Z(DIFF[20]) );
  CNR2XL U177 ( .A(A[11]), .B(n314), .Z(n311) );
  COND1X1 U178 ( .A(n203), .B(n204), .C(n187), .Z(n202) );
  CND3X1 U179 ( .A(n148), .B(n147), .C(n134), .Z(n152) );
  CND2X2 U180 ( .A(n320), .B(A[12]), .Z(n279) );
  CND2X1 U181 ( .A(A[16]), .B(n284), .Z(n229) );
  CND2XL U182 ( .A(n195), .B(n187), .Z(n40) );
  CND2IX2 U183 ( .B(n78), .A(n82), .Z(n252) );
  CANR1XL U184 ( .A(n13), .B(n37), .C(n226), .Z(n41) );
  CEOXL U185 ( .A(n42), .B(n216), .Z(DIFF[19]) );
  CANR1XL U186 ( .A(n211), .B(n110), .C(n219), .Z(n42) );
  CND2X1 U187 ( .A(n182), .B(n4), .Z(n193) );
  CND2XL U188 ( .A(n338), .B(n214), .Z(DIFF[0]) );
  COND1XL U189 ( .A(n70), .B(n71), .C(n72), .Z(n69) );
  CIVXL U190 ( .A(n73), .Z(n71) );
  CND2XL U191 ( .A(B[0]), .B(n357), .Z(n338) );
  CND2IXL U192 ( .B(B[30]), .A(A[30]), .Z(n85) );
  CNR3X1 U193 ( .A(n250), .B(n254), .C(n253), .Z(n274) );
  CND2XL U194 ( .A(n54), .B(n55), .Z(n53) );
  CNR2XL U195 ( .A(n123), .B(n179), .Z(n178) );
  CANR1XL U196 ( .A(n171), .B(n26), .C(n183), .Z(n177) );
  CND2XL U197 ( .A(n144), .B(n130), .Z(n150) );
  CND3X1 U198 ( .A(n193), .B(n192), .C(n186), .Z(n191) );
  CND2X1 U199 ( .A(n197), .B(n198), .Z(n192) );
  CND2XL U200 ( .A(n305), .B(n312), .Z(n327) );
  CND2XL U201 ( .A(n271), .B(n16), .Z(n296) );
  CND2XL U202 ( .A(n6), .B(n51), .Z(n48) );
  CND2XL U203 ( .A(n270), .B(n279), .Z(n301) );
  CND2X1 U204 ( .A(n128), .B(n129), .Z(n127) );
  CND2X1 U205 ( .A(n129), .B(n131), .Z(n125) );
  COND1XL U206 ( .A(n105), .B(n106), .C(n107), .Z(n79) );
  CND2XL U207 ( .A(n272), .B(n283), .Z(n291) );
  CND2XL U208 ( .A(n268), .B(n244), .Z(n286) );
  CENX1 U209 ( .A(n212), .B(n108), .Z(DIFF[1]) );
  CENX1 U210 ( .A(n75), .B(n76), .Z(DIFF[3]) );
  CND2XL U211 ( .A(n81), .B(n82), .Z(n75) );
  CND2X1 U212 ( .A(n77), .B(n78), .Z(n76) );
  CND2XL U213 ( .A(n79), .B(n80), .Z(n77) );
  CAN2XL U214 ( .A(n129), .B(n126), .Z(n43) );
  CENX1 U215 ( .A(n44), .B(n155), .Z(DIFF[25]) );
  CND3XL U216 ( .A(n306), .B(n305), .C(n307), .Z(n304) );
  COND1X1 U217 ( .A(n311), .B(n312), .C(n313), .Z(n303) );
  CNR2XL U218 ( .A(n308), .B(n309), .Z(n307) );
  CND2XL U219 ( .A(n147), .B(n158), .Z(n159) );
  CENXL U220 ( .A(n63), .B(n59), .Z(DIFF[6]) );
  CND2XL U221 ( .A(n7), .B(n62), .Z(n63) );
  CEOXL U222 ( .A(n45), .B(n74), .Z(DIFF[4]) );
  CAN2XL U223 ( .A(n73), .B(n72), .Z(n45) );
  CENXL U224 ( .A(n56), .B(n46), .Z(DIFF[7]) );
  CAN2XL U225 ( .A(n57), .B(n58), .Z(n46) );
  CEOXL U226 ( .A(n65), .B(n68), .Z(DIFF[5]) );
  CND2XL U227 ( .A(n67), .B(n66), .Z(n68) );
  CND2XL U228 ( .A(n213), .B(n214), .Z(n108) );
  CND2X1 U229 ( .A(n153), .B(n148), .Z(n145) );
  CNR2IX1 U230 ( .B(n268), .A(n269), .Z(n263) );
  CND3X1 U231 ( .A(n270), .B(n271), .C(n272), .Z(n269) );
  CAN2X1 U232 ( .A(n89), .B(n88), .Z(n47) );
  CND2XL U233 ( .A(n80), .B(n78), .Z(n104) );
  CND4XL U234 ( .A(n278), .B(n271), .C(n272), .D(n268), .Z(n277) );
  COND1XL U235 ( .A(n131), .B(n136), .C(n129), .Z(n135) );
  CND2XL U236 ( .A(A[0]), .B(n356), .Z(n214) );
  CND2XL U237 ( .A(A[25]), .B(n157), .Z(n143) );
  CND2XL U238 ( .A(B[26]), .B(n154), .Z(n130) );
  CND2X1 U239 ( .A(n343), .B(n214), .Z(n340) );
  CND2X1 U240 ( .A(B[1]), .B(n342), .Z(n215) );
  CND2IXL U241 ( .B(A[30]), .A(B[30]), .Z(n89) );
  CEOXL U242 ( .A(B[30]), .B(A[30]), .Z(n93) );
  CIVX1 U243 ( .A(B[20]), .Z(n206) );
  CIVX3 U244 ( .A(n271), .Z(n254) );
  CIVXL U245 ( .A(A[6]), .Z(n352) );
  CIVXL U246 ( .A(B[14]), .Z(n294) );
  CIVXL U247 ( .A(B[27]), .Z(n141) );
  CND2XL U248 ( .A(n336), .B(B[5]), .Z(n348) );
  CND2X1 U249 ( .A(B[5]), .B(n336), .Z(n67) );
  CIVX1 U250 ( .A(B[6]), .Z(n353) );
  CIVXL U251 ( .A(B[18]), .Z(n225) );
  CNR2X1 U252 ( .A(n253), .B(n254), .Z(n240) );
  CEOX1 U253 ( .A(B[31]), .B(A[31]), .Z(n83) );
  CND2X1 U254 ( .A(n199), .B(A[22]), .Z(n168) );
  CND2XL U255 ( .A(n185), .B(n168), .Z(n190) );
  CIVX2 U256 ( .A(n293), .Z(n292) );
  CENXL U257 ( .A(n301), .B(n298), .Z(DIFF[12]) );
  CEOXL U258 ( .A(n14), .B(n53), .Z(DIFF[8]) );
  CIVX2 U259 ( .A(n332), .Z(n52) );
  CND4X1 U260 ( .A(n117), .B(n125), .C(n126), .D(n127), .Z(n100) );
  CND2XL U261 ( .A(n230), .B(n229), .Z(n235) );
  CIVXL U262 ( .A(n230), .Z(n234) );
  CND2XL U263 ( .A(B[16]), .B(n285), .Z(n230) );
  CND2IXL U264 ( .B(A[17]), .A(B[17]), .Z(n221) );
  CENXL U265 ( .A(n296), .B(n293), .Z(DIFF[13]) );
  CENXL U266 ( .A(n322), .B(n323), .Z(DIFF[11]) );
  CENXL U267 ( .A(n48), .B(n21), .Z(DIFF[9]) );
  CENXL U268 ( .A(n327), .B(n325), .Z(DIFF[10]) );
  CENXL U269 ( .A(n29), .B(n235), .Z(DIFF[16]) );
  CANR1X1 U270 ( .A(n5), .B(n20), .C(n135), .Z(n133) );
  CIVX2 U271 ( .A(n62), .Z(n61) );
  CIVX2 U272 ( .A(n67), .Z(n64) );
  CENX2 U273 ( .A(n83), .B(n84), .Z(DIFF[31]) );
  CIVX2 U274 ( .A(n92), .Z(n91) );
  CND2X2 U275 ( .A(n97), .B(n88), .Z(n96) );
  CND2X2 U276 ( .A(n88), .B(n99), .Z(n95) );
  CIVX2 U277 ( .A(n100), .Z(n99) );
  CND2X2 U278 ( .A(B[29]), .B(n102), .Z(n88) );
  CIVX2 U279 ( .A(A[29]), .Z(n102) );
  CIVX2 U280 ( .A(n103), .Z(n101) );
  CND2IX1 U281 ( .B(B[29]), .A(A[29]), .Z(n92) );
  CENX1 U282 ( .A(n104), .B(n79), .Z(DIFF[2]) );
  CIVX2 U283 ( .A(n108), .Z(n106) );
  CNR2X2 U284 ( .A(n122), .B(n123), .Z(n120) );
  CIVX2 U285 ( .A(n124), .Z(n122) );
  CIVX2 U286 ( .A(n130), .Z(n128) );
  CIVX2 U287 ( .A(n132), .Z(n131) );
  CND2IX1 U288 ( .B(A[28]), .A(B[28]), .Z(n117) );
  CND2IX1 U289 ( .B(B[28]), .A(A[28]), .Z(n103) );
  CND2X2 U290 ( .A(B[27]), .B(n140), .Z(n126) );
  CIVX2 U291 ( .A(A[27]), .Z(n140) );
  CIVX2 U292 ( .A(n146), .Z(n138) );
  CND3X2 U293 ( .A(n147), .B(n148), .C(n149), .Z(n146) );
  CND2IX1 U294 ( .B(A[26]), .A(B[26]), .Z(n149) );
  CIVX2 U295 ( .A(A[26]), .Z(n154) );
  CND2IX1 U296 ( .B(B[26]), .A(A[26]), .Z(n144) );
  CND2X2 U297 ( .A(B[25]), .B(n156), .Z(n148) );
  CIVX2 U298 ( .A(A[25]), .Z(n156) );
  CIVX2 U299 ( .A(B[25]), .Z(n157) );
  CIVX2 U300 ( .A(n158), .Z(n153) );
  CIVX2 U301 ( .A(n114), .Z(n164) );
  CND2X2 U302 ( .A(n167), .B(n168), .Z(n165) );
  CND2X2 U303 ( .A(n169), .B(n119), .Z(n162) );
  CND2X2 U304 ( .A(n171), .B(n166), .Z(n170) );
  CND2X2 U305 ( .A(n172), .B(n121), .Z(n169) );
  CNR2IX2 U306 ( .B(n124), .A(n109), .Z(n172) );
  CIVX2 U307 ( .A(n173), .Z(n109) );
  CIVX2 U308 ( .A(n166), .Z(n179) );
  CND2X2 U309 ( .A(B[23]), .B(n180), .Z(n166) );
  CIVX2 U310 ( .A(A[23]), .Z(n180) );
  CIVX2 U311 ( .A(n118), .Z(n123) );
  CND2X2 U312 ( .A(A[23]), .B(n181), .Z(n118) );
  CIVX2 U313 ( .A(B[23]), .Z(n181) );
  CND3X2 U314 ( .A(n185), .B(n184), .C(n196), .Z(n167) );
  CND2X2 U315 ( .A(n186), .B(n187), .Z(n184) );
  CIVX2 U316 ( .A(n188), .Z(n171) );
  CND2X2 U317 ( .A(n189), .B(n185), .Z(n188) );
  CND2X2 U318 ( .A(n195), .B(n196), .Z(n194) );
  CND2X2 U319 ( .A(B[22]), .B(n200), .Z(n185) );
  CIVX2 U320 ( .A(A[22]), .Z(n200) );
  CND2X1 U321 ( .A(n186), .B(n197), .Z(n201) );
  CND2X2 U322 ( .A(A[21]), .B(n205), .Z(n186) );
  CIVX2 U323 ( .A(n121), .Z(n174) );
  CND2X2 U324 ( .A(n207), .B(n208), .Z(n121) );
  CND2X2 U325 ( .A(n209), .B(n210), .Z(n207) );
  CND2X2 U326 ( .A(n211), .B(n208), .Z(n173) );
  CND2X2 U327 ( .A(A[19]), .B(n217), .Z(n124) );
  CIVX2 U328 ( .A(A[19]), .Z(n218) );
  CIVX2 U329 ( .A(n223), .Z(n211) );
  CND2X2 U330 ( .A(n13), .B(n222), .Z(n223) );
  CND2X2 U331 ( .A(B[18]), .B(n224), .Z(n222) );
  CIVX2 U332 ( .A(A[18]), .Z(n224) );
  CIVX2 U333 ( .A(n220), .Z(n227) );
  CND2X2 U334 ( .A(n228), .B(n229), .Z(n220) );
  CIVX2 U335 ( .A(n252), .Z(n251) );
  CNR2X2 U336 ( .A(n257), .B(n258), .Z(n256) );
  CND2X2 U337 ( .A(n259), .B(n260), .Z(n258) );
  CNR2X2 U338 ( .A(n254), .B(n246), .Z(n259) );
  CNR2IX2 U339 ( .B(n263), .A(n264), .Z(n255) );
  CND3X2 U340 ( .A(n260), .B(n266), .C(n265), .Z(n264) );
  CIVX2 U341 ( .A(n247), .Z(n266) );
  CIVX2 U342 ( .A(n279), .Z(n278) );
  CIVX2 U343 ( .A(n283), .Z(n282) );
  CIVX2 U344 ( .A(A[16]), .Z(n285) );
  COND1X2 U345 ( .A(n254), .B(n292), .C(n16), .Z(n289) );
  COND1X2 U346 ( .A(n246), .B(n297), .C(n279), .Z(n293) );
  CIVX2 U347 ( .A(n270), .Z(n246) );
  CND2X2 U348 ( .A(B[13]), .B(n300), .Z(n271) );
  CIVX2 U349 ( .A(A[13]), .Z(n300) );
  CNR2X2 U350 ( .A(n318), .B(n308), .Z(n315) );
  CIVX2 U351 ( .A(n319), .Z(n308) );
  CIVX2 U352 ( .A(B[12]), .Z(n320) );
  CND2X2 U353 ( .A(B[12]), .B(n321), .Z(n270) );
  CIVX2 U354 ( .A(A[12]), .Z(n321) );
  CND2X2 U355 ( .A(B[11]), .B(n326), .Z(n319) );
  CIVX2 U356 ( .A(A[11]), .Z(n326) );
  COND1X2 U357 ( .A(n317), .B(n328), .C(n51), .Z(n325) );
  CIVX2 U358 ( .A(A[9]), .Z(n329) );
  CIVX2 U359 ( .A(n54), .Z(n316) );
  CND2X2 U360 ( .A(B[8]), .B(n331), .Z(n54) );
  CIVX2 U361 ( .A(A[8]), .Z(n331) );
  COND2X2 U362 ( .A(n333), .B(n334), .C(n247), .D(n70), .Z(n332) );
  CND4X2 U363 ( .A(n60), .B(n58), .C(n67), .D(n73), .Z(n247) );
  CIVX2 U364 ( .A(A[4]), .Z(n335) );
  CIVX2 U365 ( .A(n74), .Z(n70) );
  CND4X2 U366 ( .A(n252), .B(n249), .C(n81), .D(n267), .Z(n74) );
  CND3X2 U367 ( .A(n337), .B(n82), .C(n80), .Z(n267) );
  CNR2X2 U368 ( .A(n105), .B(n213), .Z(n337) );
  CIVX2 U369 ( .A(n338), .Z(n213) );
  CIVX2 U370 ( .A(n215), .Z(n105) );
  CND2X2 U371 ( .A(A[3]), .B(n339), .Z(n81) );
  CIVX2 U372 ( .A(A[2]), .Z(n341) );
  CIVX2 U373 ( .A(A[1]), .Z(n342) );
  CND2X2 U374 ( .A(B[3]), .B(n344), .Z(n82) );
  CIVX2 U375 ( .A(A[3]), .Z(n344) );
  CND2X2 U376 ( .A(A[2]), .B(n345), .Z(n78) );
  CND3X2 U377 ( .A(n346), .B(n62), .C(n57), .Z(n261) );
  CND2X2 U378 ( .A(A[7]), .B(n347), .Z(n57) );
  CND3X2 U379 ( .A(n60), .B(n348), .C(n349), .Z(n346) );
  CND2X2 U380 ( .A(n66), .B(n72), .Z(n349) );
  CND2X2 U381 ( .A(A[4]), .B(n350), .Z(n72) );
  CIVX2 U382 ( .A(B[4]), .Z(n350) );
  CND2X2 U383 ( .A(A[5]), .B(n351), .Z(n66) );
  CIVX2 U384 ( .A(B[5]), .Z(n351) );
  CND2X2 U385 ( .A(A[6]), .B(n353), .Z(n62) );
  CND2X2 U386 ( .A(B[7]), .B(n354), .Z(n58) );
  CIVX2 U387 ( .A(A[7]), .Z(n354) );
  CND2X2 U388 ( .A(B[10]), .B(n355), .Z(n305) );
  CIVX2 U389 ( .A(A[10]), .Z(n355) );
  CIVX2 U390 ( .A(B[0]), .Z(n356) );
  CIVX2 U391 ( .A(A[0]), .Z(n357) );
endmodule


module nios_2_DW01_inc_3 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181;

  CNIVXL U2 ( .A(A[13]), .Z(n1) );
  CNIVXL U3 ( .A(A[8]), .Z(n33) );
  CIVX3 U4 ( .A(n74), .Z(n70) );
  CNIVX1 U5 ( .A(A[7]), .Z(n32) );
  CNIVX4 U6 ( .A(A[1]), .Z(n2) );
  CNIVX2 U7 ( .A(A[1]), .Z(n27) );
  CIVXL U8 ( .A(A[11]), .Z(n3) );
  CIVX2 U9 ( .A(n3), .Z(n4) );
  CNR2X2 U10 ( .A(n50), .B(n51), .Z(n49) );
  CND3XL U11 ( .A(n26), .B(n29), .C(A[4]), .Z(n178) );
  CNIVX2 U12 ( .A(A[2]), .Z(n5) );
  CNIVX2 U13 ( .A(A[2]), .Z(n6) );
  CNIVX2 U14 ( .A(A[2]), .Z(n28) );
  CIVX1 U15 ( .A(n175), .Z(n17) );
  CENX1 U16 ( .A(n33), .B(n40), .Z(SUM[8]) );
  CND2X1 U17 ( .A(n41), .B(n42), .Z(n40) );
  CND2X1 U18 ( .A(n95), .B(n96), .Z(n7) );
  CND3X2 U19 ( .A(n98), .B(n97), .C(n8), .Z(n94) );
  CIVX2 U20 ( .A(n7), .Z(n8) );
  CENX1 U21 ( .A(n124), .B(n125), .Z(SUM[17]) );
  CENX1 U22 ( .A(n133), .B(n132), .Z(SUM[15]) );
  CNR2X1 U23 ( .A(n173), .B(n174), .Z(n169) );
  CND2X1 U24 ( .A(n175), .B(A[10]), .Z(n18) );
  CND2X1 U25 ( .A(A[17]), .B(A[16]), .Z(n84) );
  CND2X1 U26 ( .A(A[19]), .B(A[18]), .Z(n85) );
  CND3XL U27 ( .A(n34), .B(A[6]), .C(A[10]), .Z(n173) );
  CND2X1 U28 ( .A(n177), .B(n176), .Z(n175) );
  CENX1 U29 ( .A(n67), .B(n68), .Z(SUM[29]) );
  CENX1 U30 ( .A(A[28]), .B(n65), .Z(SUM[28]) );
  CAN2X1 U31 ( .A(n30), .B(A[4]), .Z(n9) );
  CIVX1 U32 ( .A(n30), .Z(n57) );
  CNR2X1 U33 ( .A(n144), .B(n145), .Z(n140) );
  CND2IX2 U34 ( .B(n111), .A(n112), .Z(n110) );
  CNR2X2 U35 ( .A(n113), .B(n114), .Z(n112) );
  CENX1 U36 ( .A(A[22]), .B(n92), .Z(SUM[22]) );
  CND2X1 U37 ( .A(n90), .B(n21), .Z(n92) );
  CND2XL U38 ( .A(A[7]), .B(A[6]), .Z(n145) );
  CND2X2 U39 ( .A(n29), .B(n28), .Z(n44) );
  CND2X1 U40 ( .A(A[4]), .B(n29), .Z(n118) );
  CNIVXL U41 ( .A(A[6]), .Z(n31) );
  CIVX1 U42 ( .A(n29), .Z(n61) );
  CND2X1 U43 ( .A(A[8]), .B(A[7]), .Z(n151) );
  CNIVXL U44 ( .A(A[12]), .Z(n10) );
  CND3X2 U45 ( .A(n115), .B(n116), .C(n117), .Z(n109) );
  CNR2IX1 U46 ( .B(n11), .A(n118), .Z(n38) );
  CND3X1 U47 ( .A(n37), .B(n38), .C(n36), .Z(n35) );
  CENX1 U48 ( .A(n35), .B(n34), .Z(SUM[9]) );
  CNIVX4 U49 ( .A(A[0]), .Z(n11) );
  CNIVX2 U50 ( .A(A[0]), .Z(n26) );
  CNR2X1 U51 ( .A(n151), .B(n152), .Z(n150) );
  CENX1 U52 ( .A(A[18]), .B(n123), .Z(SUM[18]) );
  CND2X1 U53 ( .A(n27), .B(n26), .Z(n43) );
  CND2XL U54 ( .A(n147), .B(n146), .Z(n14) );
  CND2X2 U55 ( .A(n12), .B(n13), .Z(n15) );
  CND2X2 U56 ( .A(n14), .B(n15), .Z(SUM[14]) );
  CIVX2 U57 ( .A(n147), .Z(n12) );
  CIVX1 U58 ( .A(n146), .Z(n13) );
  CIVXL U59 ( .A(A[14]), .Z(n147) );
  CND2X2 U60 ( .A(n17), .B(n16), .Z(n19) );
  CND2X2 U61 ( .A(n19), .B(n18), .Z(SUM[10]) );
  CIVXL U62 ( .A(A[10]), .Z(n16) );
  CNR2X1 U63 ( .A(n180), .B(n181), .Z(n176) );
  CNR2XL U64 ( .A(n77), .B(n78), .Z(n75) );
  CND2X1 U65 ( .A(n29), .B(n6), .Z(n156) );
  CND2X1 U66 ( .A(n29), .B(n5), .Z(n51) );
  CND3XL U67 ( .A(n91), .B(A[21]), .C(A[20]), .Z(n20) );
  CIVX1 U68 ( .A(n20), .Z(n21) );
  CIVX1 U69 ( .A(n93), .Z(n91) );
  CNR2IX2 U70 ( .B(A[16]), .A(n78), .Z(n124) );
  CND2X2 U71 ( .A(n54), .B(n9), .Z(n53) );
  CIVX1 U72 ( .A(n55), .Z(n54) );
  CND2X1 U73 ( .A(A[12]), .B(A[11]), .Z(n114) );
  CNR2X1 U74 ( .A(n178), .B(n179), .Z(n177) );
  CAN2XL U75 ( .A(n2), .B(n5), .Z(n115) );
  CND2XL U76 ( .A(n29), .B(n5), .Z(n143) );
  CNR2X2 U77 ( .A(n148), .B(n149), .Z(n146) );
  CND4X2 U78 ( .A(A[7]), .B(A[6]), .C(n30), .D(A[4]), .Z(n129) );
  CNR2X2 U79 ( .A(n128), .B(n129), .Z(n127) );
  CND3XL U80 ( .A(n34), .B(A[8]), .C(n30), .Z(n180) );
  CND2XL U81 ( .A(A[10]), .B(n34), .Z(n152) );
  CNIVX4 U82 ( .A(A[5]), .Z(n30) );
  CND2X1 U83 ( .A(n2), .B(n28), .Z(n59) );
  CNR2X2 U84 ( .A(n110), .B(n93), .Z(n22) );
  CNR2X4 U85 ( .A(n23), .B(n109), .Z(n107) );
  CIVX2 U86 ( .A(n22), .Z(n23) );
  CND4X1 U87 ( .A(A[19]), .B(A[18]), .C(A[17]), .D(A[16]), .Z(n93) );
  CEOX2 U88 ( .A(n162), .B(n10), .Z(SUM[12]) );
  CNR2X2 U89 ( .A(n130), .B(n131), .Z(n126) );
  CND4X1 U90 ( .A(A[11]), .B(A[10]), .C(n34), .D(A[8]), .Z(n130) );
  CND3X1 U91 ( .A(n29), .B(n30), .C(A[4]), .Z(n172) );
  CIVX1 U92 ( .A(n78), .Z(n80) );
  CENX1 U93 ( .A(A[19]), .B(n121), .Z(SUM[19]) );
  CND2X2 U94 ( .A(n127), .B(n126), .Z(n78) );
  CND2X1 U95 ( .A(A[7]), .B(A[6]), .Z(n167) );
  CND4X2 U96 ( .A(n29), .B(n6), .C(n2), .D(n11), .Z(n128) );
  CND2XL U97 ( .A(n27), .B(n11), .Z(n62) );
  CNR2X1 U98 ( .A(n143), .B(n142), .Z(n141) );
  CND2XL U99 ( .A(A[6]), .B(n30), .Z(n119) );
  CND2X1 U100 ( .A(n122), .B(A[18]), .Z(n121) );
  CAN2XL U101 ( .A(n2), .B(n6), .Z(n36) );
  CND2XL U102 ( .A(n2), .B(n5), .Z(n179) );
  CND2XL U103 ( .A(n27), .B(n11), .Z(n155) );
  CND2XL U104 ( .A(n30), .B(A[4]), .Z(n144) );
  CND2XL U105 ( .A(n2), .B(n11), .Z(n142) );
  CND2XL U106 ( .A(A[6]), .B(n30), .Z(n39) );
  CNR2X1 U107 ( .A(n101), .B(n102), .Z(n97) );
  CEOX2 U108 ( .A(A[30]), .B(n64), .Z(SUM[30]) );
  CAN2X2 U109 ( .A(n90), .B(n24), .Z(n88) );
  CAN4X1 U110 ( .A(A[21]), .B(A[22]), .C(A[20]), .D(n91), .Z(n24) );
  CND2XL U111 ( .A(n34), .B(A[8]), .Z(n138) );
  CND2IX1 U112 ( .B(n25), .A(n150), .Z(n149) );
  CND3XL U113 ( .A(A[12]), .B(A[11]), .C(A[13]), .Z(n25) );
  CNIVX4 U114 ( .A(A[3]), .Z(n29) );
  CNR2X1 U115 ( .A(n99), .B(n100), .Z(n98) );
  CNR2X1 U116 ( .A(n39), .B(n151), .Z(n37) );
  CENX1 U117 ( .A(n60), .B(n61), .Z(SUM[3]) );
  CNR2IX1 U118 ( .B(n5), .A(n62), .Z(n60) );
  CNR2X1 U119 ( .A(n155), .B(n44), .Z(n42) );
  CNR2X1 U120 ( .A(n45), .B(n46), .Z(n41) );
  CENX1 U121 ( .A(n165), .B(n6), .Z(SUM[2]) );
  CENX1 U122 ( .A(n57), .B(n56), .Z(SUM[5]) );
  CNR2X1 U123 ( .A(n119), .B(n120), .Z(n116) );
  CNR2X1 U124 ( .A(n52), .B(n57), .Z(n48) );
  CND3XL U125 ( .A(n30), .B(A[6]), .C(A[4]), .Z(n153) );
  CND2XL U126 ( .A(A[6]), .B(A[7]), .Z(n181) );
  CND2XL U127 ( .A(A[8]), .B(A[7]), .Z(n120) );
  CND2XL U128 ( .A(A[7]), .B(A[8]), .Z(n174) );
  CND2XL U129 ( .A(A[7]), .B(A[6]), .Z(n46) );
  CND2XL U130 ( .A(A[7]), .B(A[8]), .Z(n102) );
  CNR2IX1 U131 ( .B(A[28]), .A(n65), .Z(n67) );
  CND3X1 U132 ( .A(A[24]), .B(A[25]), .C(n73), .Z(n77) );
  CNR2X1 U133 ( .A(n105), .B(n106), .Z(n95) );
  CNR2X1 U134 ( .A(n65), .B(n66), .Z(n64) );
  CND2X1 U135 ( .A(A[28]), .B(A[29]), .Z(n66) );
  CEOX1 U136 ( .A(n81), .B(A[24]), .Z(SUM[24]) );
  CNR2IXL U137 ( .B(A[27]), .A(n71), .Z(n69) );
  CND3XL U138 ( .A(A[14]), .B(A[13]), .C(A[15]), .Z(n105) );
  CENX1 U139 ( .A(A[31]), .B(n63), .Z(SUM[31]) );
  CNR2X1 U140 ( .A(n103), .B(n104), .Z(n96) );
  CND3XL U141 ( .A(A[17]), .B(A[19]), .C(A[18]), .Z(n103) );
  CND3XL U142 ( .A(n34), .B(A[6]), .C(A[16]), .Z(n101) );
  CNR2X1 U143 ( .A(n138), .B(n139), .Z(n137) );
  CND2XL U144 ( .A(A[30]), .B(n64), .Z(n63) );
  CIVXL U145 ( .A(n11), .Z(SUM[0]) );
  CEOXL U146 ( .A(n2), .B(n11), .Z(SUM[1]) );
  CND3XL U147 ( .A(n5), .B(n11), .C(n2), .Z(n99) );
  CND2XL U148 ( .A(n27), .B(n26), .Z(n50) );
  CNR2IX1 U149 ( .B(n11), .A(n118), .Z(n117) );
  CND3X1 U150 ( .A(n5), .B(n11), .C(n2), .Z(n171) );
  CND3X1 U151 ( .A(n26), .B(n29), .C(A[4]), .Z(n58) );
  CND2X1 U152 ( .A(n2), .B(n11), .Z(n165) );
  CND3XL U153 ( .A(A[13]), .B(A[14]), .C(A[12]), .Z(n136) );
  CND4X1 U154 ( .A(A[15]), .B(A[14]), .C(A[13]), .D(A[12]), .Z(n131) );
  CND3XL U155 ( .A(A[14]), .B(A[15]), .C(A[13]), .Z(n111) );
  CENX2 U156 ( .A(n4), .B(n168), .Z(SUM[11]) );
  CENX1 U157 ( .A(n75), .B(n76), .Z(SUM[26]) );
  CND2IX2 U158 ( .B(n153), .A(n154), .Z(n148) );
  CND2X1 U159 ( .A(A[10]), .B(n34), .Z(n113) );
  CNIVX4 U160 ( .A(A[9]), .Z(n34) );
  CENX1 U161 ( .A(A[4]), .B(n55), .Z(SUM[4]) );
  CND3XL U162 ( .A(n29), .B(n30), .C(A[4]), .Z(n100) );
  CND2XL U163 ( .A(A[6]), .B(A[4]), .Z(n52) );
  CND2XL U164 ( .A(n30), .B(A[4]), .Z(n45) );
  CND2X1 U165 ( .A(n30), .B(A[4]), .Z(n166) );
  CNR2X1 U166 ( .A(n78), .B(n71), .Z(n81) );
  CENXL U167 ( .A(A[16]), .B(n78), .Z(SUM[16]) );
  CND2XL U168 ( .A(A[12]), .B(A[11]), .Z(n106) );
  CND2X1 U169 ( .A(A[11]), .B(A[10]), .Z(n139) );
  CND2XL U170 ( .A(A[10]), .B(A[20]), .Z(n104) );
  CND4X1 U171 ( .A(A[11]), .B(A[10]), .C(n34), .D(A[8]), .Z(n160) );
  CENX2 U172 ( .A(n32), .B(n47), .Z(SUM[7]) );
  CND2X2 U173 ( .A(n49), .B(n48), .Z(n47) );
  CENX2 U174 ( .A(n31), .B(n53), .Z(SUM[6]) );
  CNR2X2 U175 ( .A(n58), .B(n59), .Z(n56) );
  CND4X2 U176 ( .A(n29), .B(n28), .C(n27), .D(n26), .Z(n55) );
  CIVX2 U177 ( .A(A[29]), .Z(n68) );
  CND2X2 U178 ( .A(n69), .B(n70), .Z(n65) );
  CENX2 U179 ( .A(A[27]), .B(n72), .Z(SUM[27]) );
  CND2X2 U180 ( .A(n73), .B(n70), .Z(n72) );
  CND4X2 U181 ( .A(A[26]), .B(A[25]), .C(A[24]), .D(n80), .Z(n74) );
  CIVX2 U182 ( .A(A[26]), .Z(n76) );
  CIVX2 U183 ( .A(n71), .Z(n73) );
  CENX2 U184 ( .A(A[25]), .B(n79), .Z(SUM[25]) );
  CND3X2 U185 ( .A(n73), .B(n80), .C(A[24]), .Z(n79) );
  CND2X2 U186 ( .A(n82), .B(n83), .Z(n71) );
  CNR2X2 U187 ( .A(n84), .B(n85), .Z(n83) );
  CNR2X2 U188 ( .A(n86), .B(n87), .Z(n82) );
  CND2X2 U189 ( .A(A[23]), .B(A[22]), .Z(n87) );
  CND2X2 U190 ( .A(A[21]), .B(A[20]), .Z(n86) );
  CENX2 U191 ( .A(n88), .B(n89), .Z(SUM[23]) );
  CIVX2 U192 ( .A(A[23]), .Z(n89) );
  CIVX2 U193 ( .A(n78), .Z(n90) );
  CENX2 U194 ( .A(A[21]), .B(n94), .Z(SUM[21]) );
  CENX2 U195 ( .A(n108), .B(n107), .Z(SUM[20]) );
  CIVX2 U196 ( .A(A[20]), .Z(n108) );
  CIVX2 U197 ( .A(n123), .Z(n122) );
  CND3X2 U198 ( .A(A[17]), .B(A[16]), .C(n90), .Z(n123) );
  CIVX2 U199 ( .A(A[17]), .Z(n125) );
  CIVX2 U200 ( .A(A[15]), .Z(n133) );
  CNR2X2 U201 ( .A(n134), .B(n135), .Z(n132) );
  CND2IX1 U202 ( .B(n136), .A(n137), .Z(n135) );
  CND2X1 U203 ( .A(n141), .B(n140), .Z(n134) );
  CNR2X2 U204 ( .A(n165), .B(n156), .Z(n154) );
  CENX2 U205 ( .A(n1), .B(n157), .Z(SUM[13]) );
  CND3X2 U206 ( .A(n10), .B(n158), .C(n159), .Z(n157) );
  CIVX2 U207 ( .A(n160), .Z(n159) );
  CIVX2 U208 ( .A(n161), .Z(n158) );
  CNR2X2 U209 ( .A(n161), .B(n160), .Z(n162) );
  CND2X2 U210 ( .A(n164), .B(n163), .Z(n161) );
  CNR2X2 U211 ( .A(n43), .B(n44), .Z(n164) );
  CNR2X2 U212 ( .A(n166), .B(n167), .Z(n163) );
  CND2X2 U213 ( .A(n169), .B(n170), .Z(n168) );
  CNR2X2 U214 ( .A(n171), .B(n172), .Z(n170) );
endmodule


module nios_2 ( clk, rst, enable, inst_fetch, prog_count_o, data_mem_wr_o, 
        data_mem_rd_o, data_mem_addr_o, data_mem_wdata_o, data_mem_rdata_i );
  input [31:0] inst_fetch;
  output [7:0] prog_count_o;
  output [31:0] data_mem_addr_o;
  output [31:0] data_mem_wdata_o;
  input [31:0] data_mem_rdata_i;
  input clk, rst, enable;
  output data_mem_wr_o, data_mem_rd_o;
  wire   N22, N23, j_type_c, N30, N31, N32, i_type, N64, N65, N66, N67, N68,
         N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82,
         N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96,
         N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108,
         N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119,
         N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, r_type,
         N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147,
         N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158,
         N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169,
         N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180,
         N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191,
         N192, N193, N194, N195, N196, N197, N198, N199, N200, i_type_mem,
         i_type_wb_c, j_type_mem, j_type_wb_c, data_mem_rd_d, r_type_wb,
         i_type_wb, j_type_wb, \reg_mem[31][31] , \reg_mem[31][30] ,
         \reg_mem[31][29] , \reg_mem[31][28] , \reg_mem[31][27] ,
         \reg_mem[31][26] , \reg_mem[31][25] , \reg_mem[31][24] ,
         \reg_mem[31][23] , \reg_mem[31][22] , \reg_mem[31][21] ,
         \reg_mem[31][20] , \reg_mem[31][19] , \reg_mem[31][18] ,
         \reg_mem[31][17] , \reg_mem[31][16] , \reg_mem[31][15] ,
         \reg_mem[31][14] , \reg_mem[31][13] , \reg_mem[31][12] ,
         \reg_mem[31][11] , \reg_mem[31][10] , \reg_mem[31][9] ,
         \reg_mem[31][8] , \reg_mem[31][7] , \reg_mem[31][6] ,
         \reg_mem[31][5] , \reg_mem[31][4] , \reg_mem[31][3] ,
         \reg_mem[31][2] , \reg_mem[31][1] , \reg_mem[31][0] ,
         \reg_mem[30][31] , \reg_mem[30][30] , \reg_mem[30][29] ,
         \reg_mem[30][28] , \reg_mem[30][27] , \reg_mem[30][26] ,
         \reg_mem[30][25] , \reg_mem[30][24] , \reg_mem[30][23] ,
         \reg_mem[30][22] , \reg_mem[30][21] , \reg_mem[30][20] ,
         \reg_mem[30][19] , \reg_mem[30][18] , \reg_mem[30][17] ,
         \reg_mem[30][16] , \reg_mem[30][15] , \reg_mem[30][14] ,
         \reg_mem[30][13] , \reg_mem[30][12] , \reg_mem[30][11] ,
         \reg_mem[30][10] , \reg_mem[30][9] , \reg_mem[30][8] ,
         \reg_mem[30][7] , \reg_mem[30][6] , \reg_mem[30][5] ,
         \reg_mem[30][4] , \reg_mem[30][3] , \reg_mem[30][2] ,
         \reg_mem[30][1] , \reg_mem[30][0] , \reg_mem[29][31] ,
         \reg_mem[29][30] , \reg_mem[29][29] , \reg_mem[29][28] ,
         \reg_mem[29][27] , \reg_mem[29][26] , \reg_mem[29][25] ,
         \reg_mem[29][24] , \reg_mem[29][23] , \reg_mem[29][22] ,
         \reg_mem[29][21] , \reg_mem[29][20] , \reg_mem[29][19] ,
         \reg_mem[29][18] , \reg_mem[29][17] , \reg_mem[29][16] ,
         \reg_mem[29][15] , \reg_mem[29][14] , \reg_mem[29][13] ,
         \reg_mem[29][12] , \reg_mem[29][11] , \reg_mem[29][10] ,
         \reg_mem[29][9] , \reg_mem[29][8] , \reg_mem[29][7] ,
         \reg_mem[29][6] , \reg_mem[29][5] , \reg_mem[29][4] ,
         \reg_mem[29][3] , \reg_mem[29][2] , \reg_mem[29][1] ,
         \reg_mem[29][0] , \reg_mem[28][31] , \reg_mem[28][30] ,
         \reg_mem[28][29] , \reg_mem[28][28] , \reg_mem[28][27] ,
         \reg_mem[28][26] , \reg_mem[28][25] , \reg_mem[28][24] ,
         \reg_mem[28][23] , \reg_mem[28][22] , \reg_mem[28][21] ,
         \reg_mem[28][20] , \reg_mem[28][19] , \reg_mem[28][18] ,
         \reg_mem[28][17] , \reg_mem[28][16] , \reg_mem[28][15] ,
         \reg_mem[28][14] , \reg_mem[28][13] , \reg_mem[28][12] ,
         \reg_mem[28][11] , \reg_mem[28][10] , \reg_mem[28][9] ,
         \reg_mem[28][8] , \reg_mem[28][7] , \reg_mem[28][6] ,
         \reg_mem[28][5] , \reg_mem[28][4] , \reg_mem[28][3] ,
         \reg_mem[28][2] , \reg_mem[28][1] , \reg_mem[28][0] ,
         \reg_mem[27][31] , \reg_mem[27][30] , \reg_mem[27][29] ,
         \reg_mem[27][28] , \reg_mem[27][27] , \reg_mem[27][26] ,
         \reg_mem[27][25] , \reg_mem[27][24] , \reg_mem[27][23] ,
         \reg_mem[27][22] , \reg_mem[27][21] , \reg_mem[27][20] ,
         \reg_mem[27][19] , \reg_mem[27][18] , \reg_mem[27][17] ,
         \reg_mem[27][16] , \reg_mem[27][15] , \reg_mem[27][14] ,
         \reg_mem[27][13] , \reg_mem[27][12] , \reg_mem[27][11] ,
         \reg_mem[27][10] , \reg_mem[27][9] , \reg_mem[27][8] ,
         \reg_mem[27][7] , \reg_mem[27][6] , \reg_mem[27][5] ,
         \reg_mem[27][4] , \reg_mem[27][3] , \reg_mem[27][2] ,
         \reg_mem[27][1] , \reg_mem[27][0] , \reg_mem[26][31] ,
         \reg_mem[26][30] , \reg_mem[26][29] , \reg_mem[26][28] ,
         \reg_mem[26][27] , \reg_mem[26][26] , \reg_mem[26][25] ,
         \reg_mem[26][24] , \reg_mem[26][23] , \reg_mem[26][22] ,
         \reg_mem[26][21] , \reg_mem[26][20] , \reg_mem[26][19] ,
         \reg_mem[26][18] , \reg_mem[26][17] , \reg_mem[26][16] ,
         \reg_mem[26][15] , \reg_mem[26][14] , \reg_mem[26][13] ,
         \reg_mem[26][12] , \reg_mem[26][11] , \reg_mem[26][10] ,
         \reg_mem[26][9] , \reg_mem[26][8] , \reg_mem[26][7] ,
         \reg_mem[26][6] , \reg_mem[26][5] , \reg_mem[26][4] ,
         \reg_mem[26][3] , \reg_mem[26][2] , \reg_mem[26][1] ,
         \reg_mem[26][0] , \reg_mem[25][31] , \reg_mem[25][30] ,
         \reg_mem[25][29] , \reg_mem[25][28] , \reg_mem[25][27] ,
         \reg_mem[25][26] , \reg_mem[25][25] , \reg_mem[25][24] ,
         \reg_mem[25][23] , \reg_mem[25][22] , \reg_mem[25][21] ,
         \reg_mem[25][20] , \reg_mem[25][19] , \reg_mem[25][18] ,
         \reg_mem[25][17] , \reg_mem[25][16] , \reg_mem[25][15] ,
         \reg_mem[25][14] , \reg_mem[25][13] , \reg_mem[25][12] ,
         \reg_mem[25][11] , \reg_mem[25][10] , \reg_mem[25][9] ,
         \reg_mem[25][8] , \reg_mem[25][7] , \reg_mem[25][6] ,
         \reg_mem[25][5] , \reg_mem[25][4] , \reg_mem[25][3] ,
         \reg_mem[25][2] , \reg_mem[25][1] , \reg_mem[25][0] ,
         \reg_mem[24][31] , \reg_mem[24][30] , \reg_mem[24][29] ,
         \reg_mem[24][28] , \reg_mem[24][27] , \reg_mem[24][26] ,
         \reg_mem[24][25] , \reg_mem[24][24] , \reg_mem[24][23] ,
         \reg_mem[24][22] , \reg_mem[24][21] , \reg_mem[24][20] ,
         \reg_mem[24][19] , \reg_mem[24][18] , \reg_mem[24][17] ,
         \reg_mem[24][16] , \reg_mem[24][15] , \reg_mem[24][14] ,
         \reg_mem[24][13] , \reg_mem[24][12] , \reg_mem[24][11] ,
         \reg_mem[24][10] , \reg_mem[24][9] , \reg_mem[24][8] ,
         \reg_mem[24][7] , \reg_mem[24][6] , \reg_mem[24][5] ,
         \reg_mem[24][4] , \reg_mem[24][3] , \reg_mem[24][2] ,
         \reg_mem[24][1] , \reg_mem[24][0] , \reg_mem[23][31] ,
         \reg_mem[23][30] , \reg_mem[23][29] , \reg_mem[23][28] ,
         \reg_mem[23][27] , \reg_mem[23][26] , \reg_mem[23][25] ,
         \reg_mem[23][24] , \reg_mem[23][23] , \reg_mem[23][22] ,
         \reg_mem[23][21] , \reg_mem[23][20] , \reg_mem[23][19] ,
         \reg_mem[23][18] , \reg_mem[23][17] , \reg_mem[23][16] ,
         \reg_mem[23][15] , \reg_mem[23][14] , \reg_mem[23][13] ,
         \reg_mem[23][12] , \reg_mem[23][11] , \reg_mem[23][10] ,
         \reg_mem[23][9] , \reg_mem[23][8] , \reg_mem[23][7] ,
         \reg_mem[23][6] , \reg_mem[23][5] , \reg_mem[23][4] ,
         \reg_mem[23][3] , \reg_mem[23][2] , \reg_mem[23][1] ,
         \reg_mem[23][0] , \reg_mem[22][31] , \reg_mem[22][30] ,
         \reg_mem[22][29] , \reg_mem[22][28] , \reg_mem[22][27] ,
         \reg_mem[22][26] , \reg_mem[22][25] , \reg_mem[22][24] ,
         \reg_mem[22][23] , \reg_mem[22][22] , \reg_mem[22][21] ,
         \reg_mem[22][20] , \reg_mem[22][19] , \reg_mem[22][18] ,
         \reg_mem[22][17] , \reg_mem[22][16] , \reg_mem[22][15] ,
         \reg_mem[22][14] , \reg_mem[22][13] , \reg_mem[22][12] ,
         \reg_mem[22][11] , \reg_mem[22][10] , \reg_mem[22][9] ,
         \reg_mem[22][8] , \reg_mem[22][7] , \reg_mem[22][6] ,
         \reg_mem[22][5] , \reg_mem[22][4] , \reg_mem[22][3] ,
         \reg_mem[22][2] , \reg_mem[22][1] , \reg_mem[22][0] ,
         \reg_mem[21][31] , \reg_mem[21][30] , \reg_mem[21][29] ,
         \reg_mem[21][28] , \reg_mem[21][27] , \reg_mem[21][26] ,
         \reg_mem[21][25] , \reg_mem[21][24] , \reg_mem[21][23] ,
         \reg_mem[21][22] , \reg_mem[21][21] , \reg_mem[21][20] ,
         \reg_mem[21][19] , \reg_mem[21][18] , \reg_mem[21][17] ,
         \reg_mem[21][16] , \reg_mem[21][15] , \reg_mem[21][14] ,
         \reg_mem[21][13] , \reg_mem[21][12] , \reg_mem[21][11] ,
         \reg_mem[21][10] , \reg_mem[21][9] , \reg_mem[21][8] ,
         \reg_mem[21][7] , \reg_mem[21][6] , \reg_mem[21][5] ,
         \reg_mem[21][4] , \reg_mem[21][3] , \reg_mem[21][2] ,
         \reg_mem[21][1] , \reg_mem[21][0] , \reg_mem[20][31] ,
         \reg_mem[20][30] , \reg_mem[20][29] , \reg_mem[20][28] ,
         \reg_mem[20][27] , \reg_mem[20][26] , \reg_mem[20][25] ,
         \reg_mem[20][24] , \reg_mem[20][23] , \reg_mem[20][22] ,
         \reg_mem[20][21] , \reg_mem[20][20] , \reg_mem[20][19] ,
         \reg_mem[20][18] , \reg_mem[20][17] , \reg_mem[20][16] ,
         \reg_mem[20][15] , \reg_mem[20][14] , \reg_mem[20][13] ,
         \reg_mem[20][12] , \reg_mem[20][11] , \reg_mem[20][10] ,
         \reg_mem[20][9] , \reg_mem[20][8] , \reg_mem[20][7] ,
         \reg_mem[20][6] , \reg_mem[20][5] , \reg_mem[20][4] ,
         \reg_mem[20][3] , \reg_mem[20][2] , \reg_mem[20][1] ,
         \reg_mem[20][0] , \reg_mem[19][31] , \reg_mem[19][30] ,
         \reg_mem[19][29] , \reg_mem[19][28] , \reg_mem[19][27] ,
         \reg_mem[19][26] , \reg_mem[19][25] , \reg_mem[19][24] ,
         \reg_mem[19][23] , \reg_mem[19][22] , \reg_mem[19][21] ,
         \reg_mem[19][20] , \reg_mem[19][19] , \reg_mem[19][18] ,
         \reg_mem[19][17] , \reg_mem[19][16] , \reg_mem[19][15] ,
         \reg_mem[19][14] , \reg_mem[19][13] , \reg_mem[19][12] ,
         \reg_mem[19][11] , \reg_mem[19][10] , \reg_mem[19][9] ,
         \reg_mem[19][8] , \reg_mem[19][7] , \reg_mem[19][6] ,
         \reg_mem[19][5] , \reg_mem[19][4] , \reg_mem[19][3] ,
         \reg_mem[19][2] , \reg_mem[19][1] , \reg_mem[19][0] ,
         \reg_mem[18][31] , \reg_mem[18][30] , \reg_mem[18][29] ,
         \reg_mem[18][28] , \reg_mem[18][27] , \reg_mem[18][26] ,
         \reg_mem[18][25] , \reg_mem[18][24] , \reg_mem[18][23] ,
         \reg_mem[18][22] , \reg_mem[18][21] , \reg_mem[18][20] ,
         \reg_mem[18][19] , \reg_mem[18][18] , \reg_mem[18][17] ,
         \reg_mem[18][16] , \reg_mem[18][15] , \reg_mem[18][14] ,
         \reg_mem[18][13] , \reg_mem[18][12] , \reg_mem[18][11] ,
         \reg_mem[18][10] , \reg_mem[18][9] , \reg_mem[18][8] ,
         \reg_mem[18][7] , \reg_mem[18][6] , \reg_mem[18][5] ,
         \reg_mem[18][4] , \reg_mem[18][3] , \reg_mem[18][2] ,
         \reg_mem[18][1] , \reg_mem[18][0] , \reg_mem[17][31] ,
         \reg_mem[17][30] , \reg_mem[17][29] , \reg_mem[17][28] ,
         \reg_mem[17][27] , \reg_mem[17][26] , \reg_mem[17][25] ,
         \reg_mem[17][24] , \reg_mem[17][23] , \reg_mem[17][22] ,
         \reg_mem[17][21] , \reg_mem[17][20] , \reg_mem[17][19] ,
         \reg_mem[17][18] , \reg_mem[17][17] , \reg_mem[17][16] ,
         \reg_mem[17][15] , \reg_mem[17][14] , \reg_mem[17][13] ,
         \reg_mem[17][12] , \reg_mem[17][11] , \reg_mem[17][10] ,
         \reg_mem[17][9] , \reg_mem[17][8] , \reg_mem[17][7] ,
         \reg_mem[17][6] , \reg_mem[17][5] , \reg_mem[17][4] ,
         \reg_mem[17][3] , \reg_mem[17][2] , \reg_mem[17][1] ,
         \reg_mem[17][0] , \reg_mem[16][31] , \reg_mem[16][30] ,
         \reg_mem[16][29] , \reg_mem[16][28] , \reg_mem[16][27] ,
         \reg_mem[16][26] , \reg_mem[16][25] , \reg_mem[16][24] ,
         \reg_mem[16][23] , \reg_mem[16][22] , \reg_mem[16][21] ,
         \reg_mem[16][20] , \reg_mem[16][19] , \reg_mem[16][18] ,
         \reg_mem[16][17] , \reg_mem[16][16] , \reg_mem[16][15] ,
         \reg_mem[16][14] , \reg_mem[16][13] , \reg_mem[16][12] ,
         \reg_mem[16][11] , \reg_mem[16][10] , \reg_mem[16][9] ,
         \reg_mem[16][8] , \reg_mem[16][7] , \reg_mem[16][6] ,
         \reg_mem[16][5] , \reg_mem[16][4] , \reg_mem[16][3] ,
         \reg_mem[16][2] , \reg_mem[16][1] , \reg_mem[16][0] ,
         \reg_mem[15][31] , \reg_mem[15][30] , \reg_mem[15][29] ,
         \reg_mem[15][28] , \reg_mem[15][27] , \reg_mem[15][26] ,
         \reg_mem[15][25] , \reg_mem[15][24] , \reg_mem[15][23] ,
         \reg_mem[15][22] , \reg_mem[15][21] , \reg_mem[15][20] ,
         \reg_mem[15][19] , \reg_mem[15][18] , \reg_mem[15][17] ,
         \reg_mem[15][16] , \reg_mem[15][15] , \reg_mem[15][14] ,
         \reg_mem[15][13] , \reg_mem[15][12] , \reg_mem[15][11] ,
         \reg_mem[15][10] , \reg_mem[15][9] , \reg_mem[15][8] ,
         \reg_mem[15][7] , \reg_mem[15][6] , \reg_mem[15][5] ,
         \reg_mem[15][4] , \reg_mem[15][3] , \reg_mem[15][2] ,
         \reg_mem[15][1] , \reg_mem[15][0] , \reg_mem[14][31] ,
         \reg_mem[14][30] , \reg_mem[14][29] , \reg_mem[14][28] ,
         \reg_mem[14][27] , \reg_mem[14][26] , \reg_mem[14][25] ,
         \reg_mem[14][24] , \reg_mem[14][23] , \reg_mem[14][22] ,
         \reg_mem[14][21] , \reg_mem[14][20] , \reg_mem[14][19] ,
         \reg_mem[14][18] , \reg_mem[14][17] , \reg_mem[14][16] ,
         \reg_mem[14][15] , \reg_mem[14][14] , \reg_mem[14][13] ,
         \reg_mem[14][12] , \reg_mem[14][11] , \reg_mem[14][10] ,
         \reg_mem[14][9] , \reg_mem[14][8] , \reg_mem[14][7] ,
         \reg_mem[14][6] , \reg_mem[14][5] , \reg_mem[14][4] ,
         \reg_mem[14][3] , \reg_mem[14][2] , \reg_mem[14][1] ,
         \reg_mem[14][0] , \reg_mem[13][31] , \reg_mem[13][30] ,
         \reg_mem[13][29] , \reg_mem[13][28] , \reg_mem[13][27] ,
         \reg_mem[13][26] , \reg_mem[13][25] , \reg_mem[13][24] ,
         \reg_mem[13][23] , \reg_mem[13][22] , \reg_mem[13][21] ,
         \reg_mem[13][20] , \reg_mem[13][19] , \reg_mem[13][18] ,
         \reg_mem[13][17] , \reg_mem[13][16] , \reg_mem[13][15] ,
         \reg_mem[13][14] , \reg_mem[13][13] , \reg_mem[13][12] ,
         \reg_mem[13][11] , \reg_mem[13][10] , \reg_mem[13][9] ,
         \reg_mem[13][8] , \reg_mem[13][7] , \reg_mem[13][6] ,
         \reg_mem[13][5] , \reg_mem[13][4] , \reg_mem[13][3] ,
         \reg_mem[13][2] , \reg_mem[13][1] , \reg_mem[13][0] ,
         \reg_mem[12][31] , \reg_mem[12][30] , \reg_mem[12][29] ,
         \reg_mem[12][28] , \reg_mem[12][27] , \reg_mem[12][26] ,
         \reg_mem[12][25] , \reg_mem[12][24] , \reg_mem[12][23] ,
         \reg_mem[12][22] , \reg_mem[12][21] , \reg_mem[12][20] ,
         \reg_mem[12][19] , \reg_mem[12][18] , \reg_mem[12][17] ,
         \reg_mem[12][16] , \reg_mem[12][15] , \reg_mem[12][14] ,
         \reg_mem[12][13] , \reg_mem[12][12] , \reg_mem[12][11] ,
         \reg_mem[12][10] , \reg_mem[12][9] , \reg_mem[12][8] ,
         \reg_mem[12][7] , \reg_mem[12][6] , \reg_mem[12][5] ,
         \reg_mem[12][4] , \reg_mem[12][3] , \reg_mem[12][2] ,
         \reg_mem[12][1] , \reg_mem[12][0] , \reg_mem[11][31] ,
         \reg_mem[11][30] , \reg_mem[11][29] , \reg_mem[11][28] ,
         \reg_mem[11][27] , \reg_mem[11][26] , \reg_mem[11][25] ,
         \reg_mem[11][24] , \reg_mem[11][23] , \reg_mem[11][22] ,
         \reg_mem[11][21] , \reg_mem[11][20] , \reg_mem[11][19] ,
         \reg_mem[11][18] , \reg_mem[11][17] , \reg_mem[11][16] ,
         \reg_mem[11][15] , \reg_mem[11][14] , \reg_mem[11][13] ,
         \reg_mem[11][12] , \reg_mem[11][11] , \reg_mem[11][10] ,
         \reg_mem[11][9] , \reg_mem[11][8] , \reg_mem[11][7] ,
         \reg_mem[11][6] , \reg_mem[11][5] , \reg_mem[11][4] ,
         \reg_mem[11][3] , \reg_mem[11][2] , \reg_mem[11][1] ,
         \reg_mem[11][0] , \reg_mem[10][31] , \reg_mem[10][30] ,
         \reg_mem[10][29] , \reg_mem[10][28] , \reg_mem[10][27] ,
         \reg_mem[10][26] , \reg_mem[10][25] , \reg_mem[10][24] ,
         \reg_mem[10][23] , \reg_mem[10][22] , \reg_mem[10][21] ,
         \reg_mem[10][20] , \reg_mem[10][19] , \reg_mem[10][18] ,
         \reg_mem[10][17] , \reg_mem[10][16] , \reg_mem[10][15] ,
         \reg_mem[10][14] , \reg_mem[10][13] , \reg_mem[10][12] ,
         \reg_mem[10][11] , \reg_mem[10][10] , \reg_mem[10][9] ,
         \reg_mem[10][8] , \reg_mem[10][7] , \reg_mem[10][6] ,
         \reg_mem[10][5] , \reg_mem[10][4] , \reg_mem[10][3] ,
         \reg_mem[10][2] , \reg_mem[10][1] , \reg_mem[10][0] ,
         \reg_mem[9][31] , \reg_mem[9][30] , \reg_mem[9][29] ,
         \reg_mem[9][28] , \reg_mem[9][27] , \reg_mem[9][26] ,
         \reg_mem[9][25] , \reg_mem[9][24] , \reg_mem[9][23] ,
         \reg_mem[9][22] , \reg_mem[9][21] , \reg_mem[9][20] ,
         \reg_mem[9][19] , \reg_mem[9][18] , \reg_mem[9][17] ,
         \reg_mem[9][16] , \reg_mem[9][15] , \reg_mem[9][14] ,
         \reg_mem[9][13] , \reg_mem[9][12] , \reg_mem[9][11] ,
         \reg_mem[9][10] , \reg_mem[9][9] , \reg_mem[9][8] , \reg_mem[9][7] ,
         \reg_mem[9][6] , \reg_mem[9][5] , \reg_mem[9][4] , \reg_mem[9][3] ,
         \reg_mem[9][2] , \reg_mem[9][1] , \reg_mem[9][0] , \reg_mem[8][31] ,
         \reg_mem[8][30] , \reg_mem[8][29] , \reg_mem[8][28] ,
         \reg_mem[8][27] , \reg_mem[8][26] , \reg_mem[8][25] ,
         \reg_mem[8][24] , \reg_mem[8][23] , \reg_mem[8][22] ,
         \reg_mem[8][21] , \reg_mem[8][20] , \reg_mem[8][19] ,
         \reg_mem[8][18] , \reg_mem[8][17] , \reg_mem[8][16] ,
         \reg_mem[8][15] , \reg_mem[8][14] , \reg_mem[8][13] ,
         \reg_mem[8][12] , \reg_mem[8][11] , \reg_mem[8][10] , \reg_mem[8][9] ,
         \reg_mem[8][8] , \reg_mem[8][7] , \reg_mem[8][6] , \reg_mem[8][5] ,
         \reg_mem[8][4] , \reg_mem[8][3] , \reg_mem[8][2] , \reg_mem[8][1] ,
         \reg_mem[8][0] , \reg_mem[7][31] , \reg_mem[7][30] , \reg_mem[7][29] ,
         \reg_mem[7][28] , \reg_mem[7][27] , \reg_mem[7][26] ,
         \reg_mem[7][25] , \reg_mem[7][24] , \reg_mem[7][23] ,
         \reg_mem[7][22] , \reg_mem[7][21] , \reg_mem[7][20] ,
         \reg_mem[7][19] , \reg_mem[7][18] , \reg_mem[7][17] ,
         \reg_mem[7][16] , \reg_mem[7][15] , \reg_mem[7][14] ,
         \reg_mem[7][13] , \reg_mem[7][12] , \reg_mem[7][11] ,
         \reg_mem[7][10] , \reg_mem[7][9] , \reg_mem[7][8] , \reg_mem[7][7] ,
         \reg_mem[7][6] , \reg_mem[7][5] , \reg_mem[7][4] , \reg_mem[7][3] ,
         \reg_mem[7][2] , \reg_mem[7][1] , \reg_mem[7][0] , \reg_mem[6][31] ,
         \reg_mem[6][30] , \reg_mem[6][29] , \reg_mem[6][28] ,
         \reg_mem[6][27] , \reg_mem[6][26] , \reg_mem[6][25] ,
         \reg_mem[6][24] , \reg_mem[6][23] , \reg_mem[6][22] ,
         \reg_mem[6][21] , \reg_mem[6][20] , \reg_mem[6][19] ,
         \reg_mem[6][18] , \reg_mem[6][17] , \reg_mem[6][16] ,
         \reg_mem[6][15] , \reg_mem[6][14] , \reg_mem[6][13] ,
         \reg_mem[6][12] , \reg_mem[6][11] , \reg_mem[6][10] , \reg_mem[6][9] ,
         \reg_mem[6][8] , \reg_mem[6][7] , \reg_mem[6][6] , \reg_mem[6][5] ,
         \reg_mem[6][4] , \reg_mem[6][3] , \reg_mem[6][2] , \reg_mem[6][1] ,
         \reg_mem[6][0] , \reg_mem[5][31] , \reg_mem[5][30] , \reg_mem[5][29] ,
         \reg_mem[5][28] , \reg_mem[5][27] , \reg_mem[5][26] ,
         \reg_mem[5][25] , \reg_mem[5][24] , \reg_mem[5][23] ,
         \reg_mem[5][22] , \reg_mem[5][21] , \reg_mem[5][20] ,
         \reg_mem[5][19] , \reg_mem[5][18] , \reg_mem[5][17] ,
         \reg_mem[5][16] , \reg_mem[5][15] , \reg_mem[5][14] ,
         \reg_mem[5][13] , \reg_mem[5][12] , \reg_mem[5][11] ,
         \reg_mem[5][10] , \reg_mem[5][9] , \reg_mem[5][8] , \reg_mem[5][7] ,
         \reg_mem[5][6] , \reg_mem[5][5] , \reg_mem[5][4] , \reg_mem[5][3] ,
         \reg_mem[5][2] , \reg_mem[5][1] , \reg_mem[5][0] , \reg_mem[4][31] ,
         \reg_mem[4][30] , \reg_mem[4][29] , \reg_mem[4][28] ,
         \reg_mem[4][27] , \reg_mem[4][26] , \reg_mem[4][25] ,
         \reg_mem[4][24] , \reg_mem[4][23] , \reg_mem[4][22] ,
         \reg_mem[4][21] , \reg_mem[4][20] , \reg_mem[4][19] ,
         \reg_mem[4][18] , \reg_mem[4][17] , \reg_mem[4][16] ,
         \reg_mem[4][15] , \reg_mem[4][14] , \reg_mem[4][13] ,
         \reg_mem[4][12] , \reg_mem[4][11] , \reg_mem[4][10] , \reg_mem[4][9] ,
         \reg_mem[4][8] , \reg_mem[4][7] , \reg_mem[4][6] , \reg_mem[4][5] ,
         \reg_mem[4][4] , \reg_mem[4][3] , \reg_mem[4][2] , \reg_mem[4][1] ,
         \reg_mem[4][0] , \reg_mem[3][31] , \reg_mem[3][30] , \reg_mem[3][29] ,
         \reg_mem[3][28] , \reg_mem[3][27] , \reg_mem[3][26] ,
         \reg_mem[3][25] , \reg_mem[3][24] , \reg_mem[3][23] ,
         \reg_mem[3][22] , \reg_mem[3][21] , \reg_mem[3][20] ,
         \reg_mem[3][19] , \reg_mem[3][18] , \reg_mem[3][17] ,
         \reg_mem[3][16] , \reg_mem[3][15] , \reg_mem[3][14] ,
         \reg_mem[3][13] , \reg_mem[3][12] , \reg_mem[3][11] ,
         \reg_mem[3][10] , \reg_mem[3][9] , \reg_mem[3][8] , \reg_mem[3][7] ,
         \reg_mem[3][6] , \reg_mem[3][5] , \reg_mem[3][4] , \reg_mem[3][3] ,
         \reg_mem[3][2] , \reg_mem[3][1] , \reg_mem[3][0] , \reg_mem[2][31] ,
         \reg_mem[2][30] , \reg_mem[2][29] , \reg_mem[2][28] ,
         \reg_mem[2][27] , \reg_mem[2][26] , \reg_mem[2][25] ,
         \reg_mem[2][24] , \reg_mem[2][23] , \reg_mem[2][22] ,
         \reg_mem[2][21] , \reg_mem[2][20] , \reg_mem[2][19] ,
         \reg_mem[2][18] , \reg_mem[2][17] , \reg_mem[2][16] ,
         \reg_mem[2][15] , \reg_mem[2][14] , \reg_mem[2][13] ,
         \reg_mem[2][12] , \reg_mem[2][11] , \reg_mem[2][10] , \reg_mem[2][9] ,
         \reg_mem[2][8] , \reg_mem[2][7] , \reg_mem[2][6] , \reg_mem[2][5] ,
         \reg_mem[2][4] , \reg_mem[2][3] , \reg_mem[2][2] , \reg_mem[2][1] ,
         \reg_mem[2][0] , \reg_mem[1][31] , \reg_mem[1][30] , \reg_mem[1][29] ,
         \reg_mem[1][28] , \reg_mem[1][27] , \reg_mem[1][26] ,
         \reg_mem[1][25] , \reg_mem[1][24] , \reg_mem[1][23] ,
         \reg_mem[1][22] , \reg_mem[1][21] , \reg_mem[1][20] ,
         \reg_mem[1][19] , \reg_mem[1][18] , \reg_mem[1][17] ,
         \reg_mem[1][16] , \reg_mem[1][15] , \reg_mem[1][14] ,
         \reg_mem[1][13] , \reg_mem[1][12] , \reg_mem[1][11] ,
         \reg_mem[1][10] , \reg_mem[1][9] , \reg_mem[1][8] , \reg_mem[1][7] ,
         \reg_mem[1][6] , \reg_mem[1][5] , \reg_mem[1][4] , \reg_mem[1][3] ,
         \reg_mem[1][2] , \reg_mem[1][1] , \reg_mem[1][0] , \reg_mem[0][31] ,
         \reg_mem[0][30] , \reg_mem[0][29] , \reg_mem[0][28] ,
         \reg_mem[0][27] , \reg_mem[0][26] , \reg_mem[0][25] ,
         \reg_mem[0][24] , \reg_mem[0][23] , \reg_mem[0][22] ,
         \reg_mem[0][21] , \reg_mem[0][20] , \reg_mem[0][19] ,
         \reg_mem[0][18] , \reg_mem[0][17] , \reg_mem[0][16] ,
         \reg_mem[0][15] , \reg_mem[0][14] , \reg_mem[0][13] ,
         \reg_mem[0][12] , \reg_mem[0][11] , \reg_mem[0][10] , \reg_mem[0][9] ,
         \reg_mem[0][8] , \reg_mem[0][7] , \reg_mem[0][6] , \reg_mem[0][5] ,
         \reg_mem[0][4] , \reg_mem[0][3] , \reg_mem[0][2] , \reg_mem[0][1] ,
         \reg_mem[0][0] , N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N232, r_type_mem, j_type, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, n98, n99, n100, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n248, n249, n338, n339, n340, n341, n342, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, \twos_comp[9] , \twos_comp[8] ,
         \twos_comp[7] , \twos_comp[6] , \twos_comp[5] , \twos_comp[4] ,
         \twos_comp[3] , \twos_comp[31] , \twos_comp[30] , \twos_comp[2] ,
         \twos_comp[29] , \twos_comp[28] , \twos_comp[27] , \twos_comp[26] ,
         \twos_comp[25] , \twos_comp[24] , \twos_comp[23] , \twos_comp[22] ,
         \twos_comp[21] , \twos_comp[20] , \twos_comp[1] , \twos_comp[19] ,
         \twos_comp[18] , \twos_comp[17] , \twos_comp[16] , \twos_comp[15] ,
         \twos_comp[14] , \twos_comp[13] , \twos_comp[12] , \twos_comp[11] ,
         \twos_comp[10] , \twos_comp[0] , \dp_cluster_0/N63 ,
         \dp_cluster_0/N62 , \dp_cluster_0/N61 , \dp_cluster_0/N60 ,
         \dp_cluster_0/N58 , \dp_cluster_0/N57 , \dp_cluster_0/N56 ,
         \dp_cluster_0/N55 , \dp_cluster_0/N54 , \dp_cluster_0/N52 ,
         \dp_cluster_0/N51 , \dp_cluster_0/N50 , \dp_cluster_0/N49 ,
         \dp_cluster_0/N48 , \dp_cluster_0/N47 , \dp_cluster_0/N46 ,
         \dp_cluster_0/N45 , \dp_cluster_0/N44 , \dp_cluster_0/N43 ,
         \dp_cluster_0/N42 , \dp_cluster_0/N41 , \dp_cluster_0/N40 ,
         \dp_cluster_0/N39 , \dp_cluster_0/N38 , \dp_cluster_0/N37 ,
         \dp_cluster_0/N36 , \dp_cluster_0/N35 , \dp_cluster_0/N34 ,
         \dp_cluster_0/N33 , net15031, net76653, net76768, net76776, net76777,
         net76796, net77918, net77950, net78042, net78074, net78097, net78475,
         net78478, net78495, net78497, net78498, net78599, net78602, net78619,
         net78621, net78622, net78726, net78759, net78790, net78792, net78793,
         net78797, net79032, net79033, net79122, net79123, net79406, net79407,
         net79408, net79409, net79475, net79476, net79481, net79482, net79756,
         net79770, net80177, net80178, net81923, net81919, net81917, net81907,
         net81905, net81901, net81971, net81959, net81957, net81951, net81947,
         net81945, net81941, net82011, net81999, net81997, net81991, net81987,
         net81985, net81981, net82051, net82043, net82039, net82037, net82031,
         net82027, net82025, net82021, net82403, net82399, net82387, net82385,
         net82381, net82379, net82377, net82443, net82439, net82437, net82427,
         net82425, net82421, net82491, net82489, net82485, net82483, net82479,
         net82477, net82473, net82469, net82465, net82463, net82461, net82459,
         net82457, net82533, net82529, net82527, net82523, net82521, net82519,
         net82517, net82515, net82513, net82509, net82507, net82505, net82503,
         net82501, net82499, net82497, net82571, net82557, net82549, net82543,
         net82541, net82539, net82537, net82611, net82609, net82605, net82603,
         net82599, net82597, net82593, net82591, net82587, net82585, net82583,
         net82581, net82579, net82577, net82643, net82639, net82627, net82625,
         net82621, net82619, net82617, net82689, net82683, net82679, net82677,
         net82667, net82665, net82869, net82867, net82865, net82863, net82861,
         net82859, net83055, net83054, net83059, net83058, net83073, net83072,
         net83077, net83076, net83575, net83592, net86657, net86659, net86675,
         net86939, net86999, net87043, net87042, net87281, net87280, net87279,
         net87278, net87277, net87276, net87275, net87273, net87272, net87271,
         net87269, net87268, net87267, net87266, net87265, net87263, net87262,
         net87261, net87260, net87258, net87256, net87255, net87253, net87252,
         net87251, net87250, net87248, net87247, net87243, net87242, net87241,
         net87239, net87238, net87237, net87236, net87235, net87234, net87233,
         net87231, net87230, net87412, net87411, net87410, net87409, net87408,
         net87407, net87406, net87405, net87404, net87403, net87402, net87401,
         net87400, net87399, net87398, net87397, net87396, net87395, net87394,
         net87393, net87392, net87391, net87389, net87388, net87387, net87386,
         net87385, net87380, net87379, net87378, net87377, net87376, net87374,
         net87372, net87368, net87483, net87489, net87488, net87545, net87544,
         net87542, net87541, net87540, net87538, net87537, net87533, net87532,
         net87531, net87530, net87529, net87526, net87525, net87524, net87523,
         net87522, net87521, net87520, net87519, net87518, net87516, net87514,
         net87513, net87512, net87511, net87510, net87508, net87507, net87642,
         net87640, net87639, net87638, net87637, net87636, net87635, net87634,
         net87633, net87632, net87631, net87630, net87629, net87628, net87627,
         net87626, net87625, net87624, net87623, net87619, net87691, net87730,
         net87728, net87727, net87725, net87724, net87723, net87722, net87720,
         net87719, net87718, net87717, net87716, net87715, net87714, net87710,
         net87709, net87708, net87706, net87705, net87704, net87703, net87702,
         net87701, net87699, net87698, net87697, net87782, net87809, net87807,
         net87806, net87804, net87803, net87802, net87800, net87799, net87798,
         net87797, net87795, net87794, net87793, net87791, net87790, net87789,
         net87856, net87863, net87990, net88101, net88116, net88115, net88155,
         net88166, net87836, net87835, net87781, net78798, net78795, net78496,
         net86647, net80186, net80185, net80176, net80175, net76798, net78502,
         net78494, net78493, net78477, net78476, net78620, net87618, net78626,
         net78618, net78617, net78601, net78600, net87620, net78098, net87700,
         net87622, net78090, net78089, net78073, net78041, net87788, net77970,
         net77969, net77967, net88175, net87786, net77974, net77966, net77965,
         net77949, net77917, net87787, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1692, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1848, n1849, n1851, n1852, n1854, n1855, n1857, n1858, n1860, n1861,
         n1863, n1864, n1866, n1867, n1869, n1870, n1872, n1873, n1875, n1876,
         n1877, n1879, n1880, n1881, n1883, n1884, n1886, n1887, n1889, n1890,
         n1891, n1892, n1894, n1895, n1896, n1898, n1899, n1901, n1902, n1904,
         n1905, n1907, n1908, n1910, n1911, n1913, n1915, n1917, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1927, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268;
  wire   [31:0] regA;
  wire   [31:0] immi_val;
  wire   [31:0] alu_op_c;
  wire   [7:0] prog_count_c;
  wire   [4:0] regc_addr_c;
  wire   [31:0] immi_val_c;
  wire   [10:0] opcode_ext_c;
  wire   [5:0] opcode_ex;
  wire   [10:0] opcode_ext_ex;
  wire   [31:0] regB;
  wire   [7:0] prog_count_ex;
  wire   [5:0] opcode_mem;
  wire   [31:0] alu_op;
  wire   [31:0] regB_mem;
  wire   [31:0] alu_op_wb;
  wire   [4:0] regb_addr_wb;
  wire   [4:0] regc_addr_wb;
  wire   [4:0] regb_addr;
  wire   [4:0] regc_addr;
  wire   [4:0] regc_addr_mem;
  wire   [4:0] regb_addr_mem;
  wire   [7:0] prog_count_de;
  assign prog_count_o[0] = N22;
  assign prog_count_o[1] = N23;

  CFD2X1 \immi_val_reg[26]  ( .D(n5237), .CP(clk), .CD(rst), .Q(immi_val[26]), 
        .QN(\dp_cluster_0/N37 ) );
  CFD2X1 \immi_val_reg[23]  ( .D(immi_val_c[23]), .CP(clk), .CD(rst), .Q(
        immi_val[23]), .QN(\dp_cluster_0/N40 ) );
  CFD2X1 \immi_val_reg[22]  ( .D(immi_val_c[22]), .CP(clk), .CD(rst), .Q(
        immi_val[22]), .QN(\dp_cluster_0/N41 ) );
  CFD2X1 \immi_val_reg[21]  ( .D(immi_val_c[21]), .CP(clk), .CD(rst), .Q(
        immi_val[21]), .QN(\dp_cluster_0/N42 ) );
  CFD2X1 \immi_val_reg[20]  ( .D(immi_val_c[20]), .CP(clk), .CD(rst), .Q(
        immi_val[20]), .QN(\dp_cluster_0/N43 ) );
  CFD2X1 \immi_val_reg[19]  ( .D(immi_val_c[19]), .CP(clk), .CD(rst), .Q(
        immi_val[19]), .QN(\dp_cluster_0/N44 ) );
  CFD2X1 \immi_val_reg[17]  ( .D(immi_val_c[17]), .CP(clk), .CD(rst), .Q(
        immi_val[17]), .QN(\dp_cluster_0/N46 ) );
  CFD2X1 \immi_val_reg[16]  ( .D(immi_val_c[16]), .CP(clk), .CD(rst), .Q(
        immi_val[16]), .QN(\dp_cluster_0/N47 ) );
  CFD2X1 \immi_val_reg[15]  ( .D(immi_val_c[15]), .CP(clk), .CD(rst), .Q(
        immi_val[15]), .QN(\dp_cluster_0/N48 ) );
  CFD2X1 \immi_val_reg[14]  ( .D(immi_val_c[14]), .CP(clk), .CD(rst), .Q(
        immi_val[14]), .QN(\dp_cluster_0/N49 ) );
  CFD2X1 \immi_val_reg[13]  ( .D(immi_val_c[13]), .CP(clk), .CD(rst), .Q(
        immi_val[13]), .QN(\dp_cluster_0/N50 ) );
  CFD2X1 \immi_val_reg[12]  ( .D(immi_val_c[12]), .CP(clk), .CD(rst), .Q(
        immi_val[12]), .QN(\dp_cluster_0/N51 ) );
  CFD2X1 \immi_val_reg[11]  ( .D(immi_val_c[11]), .CP(clk), .CD(rst), .Q(
        immi_val[11]), .QN(\dp_cluster_0/N52 ) );
  CFD2X1 \immi_val_reg[9]  ( .D(immi_val_c[9]), .CP(clk), .CD(rst), .Q(
        immi_val[9]), .QN(\dp_cluster_0/N54 ) );
  CFD2X1 \immi_val_reg[8]  ( .D(immi_val_c[8]), .CP(clk), .CD(rst), .Q(
        immi_val[8]), .QN(\dp_cluster_0/N55 ) );
  CFD2X1 \immi_val_reg[7]  ( .D(immi_val_c[7]), .CP(clk), .CD(rst), .Q(
        immi_val[7]), .QN(\dp_cluster_0/N56 ) );
  CFD2X1 \immi_val_reg[6]  ( .D(immi_val_c[6]), .CP(clk), .CD(rst), .Q(
        immi_val[6]), .QN(\dp_cluster_0/N57 ) );
  CFD2X1 \immi_val_reg[5]  ( .D(immi_val_c[5]), .CP(clk), .CD(rst), .Q(
        immi_val[5]), .QN(\dp_cluster_0/N58 ) );
  CFD2X1 \immi_val_reg[3]  ( .D(immi_val_c[3]), .CP(clk), .CD(rst), .Q(
        immi_val[3]), .QN(\dp_cluster_0/N60 ) );
  CFD2X1 \immi_val_reg[2]  ( .D(immi_val_c[2]), .CP(clk), .CD(rst), .Q(
        immi_val[2]), .QN(\dp_cluster_0/N61 ) );
  CFD2X1 \immi_val_reg[1]  ( .D(immi_val_c[1]), .CP(clk), .CD(rst), .Q(
        immi_val[1]), .QN(\dp_cluster_0/N62 ) );
  CFD2X1 \immi_val_reg[0]  ( .D(immi_val_c[0]), .CP(clk), .CD(rst), .Q(
        immi_val[0]), .QN(\dp_cluster_0/N63 ) );
  CNR2X2 U75 ( .A(n5265), .B(n207), .Z(n210) );
  CAN3X2 U94 ( .A(n5266), .B(n5267), .C(n230), .Z(n200) );
  CAN3X2 U96 ( .A(n229), .B(n5266), .C(n230), .Z(n202) );
  CAN3X2 U98 ( .A(n231), .B(n5267), .C(n230), .Z(n204) );
  CNR2IX2 U100 ( .B(n207), .A(n5265), .Z(n228) );
  CAN3X2 U103 ( .A(n231), .B(n229), .C(n230), .Z(n206) );
  CANR2X2 U106 ( .A(regc_addr_wb[1]), .B(n240), .C(regb_addr_wb[1]), .D(n2117), 
        .Z(n231) );
  CAN3X2 U109 ( .A(n243), .B(n5268), .C(j_type_mem), .Z(j_type_wb_c) );
  CAOR2X1 U422 ( .A(\reg_mem[31][31] ), .B(n2434), .C(n2438), .D(n2269), .Z(
        n352) );
  CAOR2X1 U423 ( .A(\reg_mem[31][30] ), .B(n2434), .C(n2436), .D(n2267), .Z(
        n353) );
  CAOR2X1 U424 ( .A(\reg_mem[31][29] ), .B(n2434), .C(n2437), .D(n2265), .Z(
        n354) );
  CAOR2X1 U425 ( .A(\reg_mem[31][28] ), .B(n2434), .C(n2436), .D(n2263), .Z(
        n355) );
  CAOR2X1 U426 ( .A(\reg_mem[31][27] ), .B(n2434), .C(n2438), .D(n2261), .Z(
        n356) );
  CAOR2X1 U427 ( .A(\reg_mem[31][26] ), .B(n2434), .C(n2437), .D(n2259), .Z(
        n357) );
  CAOR2X1 U428 ( .A(\reg_mem[31][25] ), .B(n2434), .C(n2438), .D(n2257), .Z(
        n358) );
  CAOR2X1 U429 ( .A(\reg_mem[31][24] ), .B(n2434), .C(n2438), .D(n2255), .Z(
        n359) );
  CAOR2X1 U430 ( .A(\reg_mem[31][23] ), .B(n2433), .C(n2437), .D(n2253), .Z(
        n360) );
  CAOR2X1 U431 ( .A(\reg_mem[31][22] ), .B(n2433), .C(n2436), .D(n2251), .Z(
        n361) );
  CAOR2X1 U432 ( .A(\reg_mem[31][21] ), .B(n2433), .C(n2438), .D(n2249), .Z(
        n362) );
  CAOR2X1 U433 ( .A(\reg_mem[31][20] ), .B(n2433), .C(n2438), .D(n2247), .Z(
        n363) );
  CAOR2X1 U434 ( .A(\reg_mem[31][19] ), .B(n2433), .C(n2437), .D(n2245), .Z(
        n364) );
  CAOR2X1 U435 ( .A(\reg_mem[31][18] ), .B(n2433), .C(n2436), .D(n2243), .Z(
        n365) );
  CAOR2X1 U436 ( .A(\reg_mem[31][17] ), .B(n2433), .C(n2437), .D(n2241), .Z(
        n366) );
  CAOR2X1 U437 ( .A(\reg_mem[31][16] ), .B(n2433), .C(n2437), .D(n2239), .Z(
        n367) );
  CAOR2X1 U438 ( .A(\reg_mem[31][15] ), .B(n2433), .C(n2436), .D(n2237), .Z(
        n368) );
  CAOR2X1 U439 ( .A(\reg_mem[31][14] ), .B(n2433), .C(n2436), .D(n2235), .Z(
        n369) );
  CAOR2X1 U440 ( .A(\reg_mem[31][13] ), .B(n2433), .C(n2435), .D(net83055), 
        .Z(n370) );
  CAOR2X1 U441 ( .A(\reg_mem[31][12] ), .B(n2433), .C(n2437), .D(n2233), .Z(
        n371) );
  CAOR2X1 U442 ( .A(\reg_mem[31][11] ), .B(n2432), .C(n2435), .D(net83059), 
        .Z(n372) );
  CAOR2X1 U443 ( .A(\reg_mem[31][10] ), .B(n2432), .C(n2437), .D(n2231), .Z(
        n373) );
  CAOR2X1 U444 ( .A(\reg_mem[31][9] ), .B(n2432), .C(n2435), .D(n2229), .Z(
        n374) );
  CAOR2X1 U445 ( .A(\reg_mem[31][8] ), .B(n2432), .C(n2437), .D(n2227), .Z(
        n375) );
  CAOR2X1 U446 ( .A(\reg_mem[31][7] ), .B(n2432), .C(n2437), .D(n2225), .Z(
        n376) );
  CAOR2X1 U447 ( .A(\reg_mem[31][6] ), .B(n2432), .C(n2435), .D(n2223), .Z(
        n377) );
  CAOR2X1 U448 ( .A(\reg_mem[31][5] ), .B(n2432), .C(n2437), .D(n2221), .Z(
        n378) );
  CAOR2X1 U449 ( .A(\reg_mem[31][4] ), .B(n2432), .C(n2437), .D(net83073), .Z(
        n379) );
  CAOR2X1 U450 ( .A(\reg_mem[31][3] ), .B(n2432), .C(n2435), .D(n2219), .Z(
        n380) );
  CAOR2X1 U451 ( .A(\reg_mem[31][2] ), .B(n2432), .C(n2435), .D(net83077), .Z(
        n381) );
  CAOR2X1 U452 ( .A(\reg_mem[31][1] ), .B(n2432), .C(n2438), .D(n2217), .Z(
        n382) );
  CAOR2X1 U453 ( .A(\reg_mem[31][0] ), .B(n2432), .C(n2437), .D(n2215), .Z(
        n383) );
  CAOR2X1 U454 ( .A(\reg_mem[30][31] ), .B(n2427), .C(n2431), .D(n2268), .Z(
        n384) );
  CAOR2X1 U455 ( .A(\reg_mem[30][30] ), .B(n2427), .C(n2430), .D(n2266), .Z(
        n385) );
  CAOR2X1 U456 ( .A(\reg_mem[30][29] ), .B(n2427), .C(n2430), .D(n2264), .Z(
        n386) );
  CAOR2X1 U457 ( .A(\reg_mem[30][28] ), .B(n2427), .C(n2430), .D(n2262), .Z(
        n387) );
  CAOR2X1 U458 ( .A(\reg_mem[30][27] ), .B(n2427), .C(n2431), .D(n2260), .Z(
        n388) );
  CAOR2X1 U459 ( .A(\reg_mem[30][26] ), .B(n2427), .C(n2430), .D(n2258), .Z(
        n389) );
  CAOR2X1 U460 ( .A(\reg_mem[30][25] ), .B(n2427), .C(n2431), .D(n2256), .Z(
        n390) );
  CAOR2X1 U461 ( .A(\reg_mem[30][24] ), .B(n2427), .C(n2431), .D(n2254), .Z(
        n391) );
  CAOR2X1 U462 ( .A(\reg_mem[30][23] ), .B(n2426), .C(n2430), .D(n2252), .Z(
        n392) );
  CAOR2X1 U463 ( .A(\reg_mem[30][22] ), .B(n2426), .C(n2430), .D(n2250), .Z(
        n393) );
  CAOR2X1 U464 ( .A(\reg_mem[30][21] ), .B(n2426), .C(n2431), .D(n2248), .Z(
        n394) );
  CAOR2X1 U465 ( .A(\reg_mem[30][20] ), .B(n2426), .C(n2431), .D(n2246), .Z(
        n395) );
  CAOR2X1 U466 ( .A(\reg_mem[30][19] ), .B(n2426), .C(n2430), .D(n2244), .Z(
        n396) );
  CAOR2X1 U467 ( .A(\reg_mem[30][18] ), .B(n2426), .C(n2430), .D(n2242), .Z(
        n397) );
  CAOR2X1 U468 ( .A(\reg_mem[30][17] ), .B(n2426), .C(n2430), .D(n2240), .Z(
        n398) );
  CAOR2X1 U469 ( .A(\reg_mem[30][16] ), .B(n2426), .C(n2430), .D(n2238), .Z(
        n399) );
  CAOR2X1 U470 ( .A(\reg_mem[30][15] ), .B(n2426), .C(n2430), .D(n2236), .Z(
        n400) );
  CAOR2X1 U471 ( .A(\reg_mem[30][14] ), .B(n2426), .C(n2430), .D(n2234), .Z(
        n401) );
  CAOR2X1 U472 ( .A(\reg_mem[30][13] ), .B(n2426), .C(n2429), .D(net83054), 
        .Z(n402) );
  CAOR2X1 U473 ( .A(\reg_mem[30][12] ), .B(n2426), .C(n2428), .D(n2232), .Z(
        n403) );
  CAOR2X1 U474 ( .A(\reg_mem[30][11] ), .B(n2425), .C(n2429), .D(net83058), 
        .Z(n404) );
  CAOR2X1 U475 ( .A(\reg_mem[30][10] ), .B(n2425), .C(n2428), .D(n2230), .Z(
        n405) );
  CAOR2X1 U476 ( .A(\reg_mem[30][9] ), .B(n2425), .C(n2429), .D(n2228), .Z(
        n406) );
  CAOR2X1 U477 ( .A(\reg_mem[30][8] ), .B(n2425), .C(n2428), .D(n2226), .Z(
        n407) );
  CAOR2X1 U478 ( .A(\reg_mem[30][7] ), .B(n2425), .C(n2429), .D(n2224), .Z(
        n408) );
  CAOR2X1 U479 ( .A(\reg_mem[30][6] ), .B(n2425), .C(n2428), .D(n2222), .Z(
        n409) );
  CAOR2X1 U480 ( .A(\reg_mem[30][5] ), .B(n2425), .C(n2429), .D(n2220), .Z(
        n410) );
  CAOR2X1 U481 ( .A(\reg_mem[30][4] ), .B(n2425), .C(n2429), .D(net83072), .Z(
        n411) );
  CAOR2X1 U482 ( .A(\reg_mem[30][3] ), .B(n2425), .C(n2428), .D(n2218), .Z(
        n412) );
  CAOR2X1 U483 ( .A(\reg_mem[30][2] ), .B(n2425), .C(n2428), .D(net83076), .Z(
        n413) );
  CAOR2X1 U484 ( .A(\reg_mem[30][1] ), .B(n2425), .C(n2431), .D(n2216), .Z(
        n414) );
  CAOR2X1 U485 ( .A(\reg_mem[30][0] ), .B(n2425), .C(n2430), .D(n2214), .Z(
        n415) );
  CAOR2X1 U486 ( .A(\reg_mem[29][31] ), .B(n2420), .C(n2422), .D(n159), .Z(
        n416) );
  CAOR2X1 U487 ( .A(\reg_mem[29][30] ), .B(n2420), .C(n2421), .D(n160), .Z(
        n417) );
  CAOR2X1 U488 ( .A(\reg_mem[29][29] ), .B(n2420), .C(n2424), .D(n161), .Z(
        n418) );
  CAOR2X1 U489 ( .A(\reg_mem[29][28] ), .B(n2420), .C(n2423), .D(n162), .Z(
        n419) );
  CAOR2X1 U490 ( .A(\reg_mem[29][27] ), .B(n2420), .C(n2423), .D(n163), .Z(
        n420) );
  CAOR2X1 U491 ( .A(\reg_mem[29][26] ), .B(n2420), .C(n2422), .D(n164), .Z(
        n421) );
  CAOR2X1 U492 ( .A(\reg_mem[29][25] ), .B(n2420), .C(n2422), .D(n165), .Z(
        n422) );
  CAOR2X1 U493 ( .A(\reg_mem[29][24] ), .B(n2420), .C(n2422), .D(n166), .Z(
        n423) );
  CAOR2X1 U494 ( .A(\reg_mem[29][23] ), .B(n2419), .C(n2424), .D(n167), .Z(
        n424) );
  CAOR2X1 U495 ( .A(\reg_mem[29][22] ), .B(n2419), .C(n2423), .D(n168), .Z(
        n425) );
  CAOR2X1 U496 ( .A(\reg_mem[29][21] ), .B(n2419), .C(n2422), .D(n169), .Z(
        n426) );
  CAOR2X1 U497 ( .A(\reg_mem[29][20] ), .B(n2419), .C(n2422), .D(n170), .Z(
        n427) );
  CAOR2X1 U498 ( .A(\reg_mem[29][19] ), .B(n2419), .C(n2424), .D(n171), .Z(
        n428) );
  CAOR2X1 U499 ( .A(\reg_mem[29][18] ), .B(n2419), .C(n2423), .D(n172), .Z(
        n429) );
  CAOR2X1 U500 ( .A(\reg_mem[29][17] ), .B(n2419), .C(n2424), .D(n173), .Z(
        n430) );
  CAOR2X1 U501 ( .A(\reg_mem[29][16] ), .B(n2419), .C(n2424), .D(n174), .Z(
        n431) );
  CAOR2X1 U502 ( .A(\reg_mem[29][15] ), .B(n2419), .C(n2423), .D(n175), .Z(
        n432) );
  CAOR2X1 U503 ( .A(\reg_mem[29][14] ), .B(n2419), .C(n2423), .D(n176), .Z(
        n433) );
  CAOR2X1 U504 ( .A(\reg_mem[29][13] ), .B(n2419), .C(n2422), .D(n177), .Z(
        n434) );
  CAOR2X1 U505 ( .A(\reg_mem[29][12] ), .B(n2419), .C(n2421), .D(n178), .Z(
        n435) );
  CAOR2X1 U506 ( .A(\reg_mem[29][11] ), .B(n2418), .C(n2422), .D(n179), .Z(
        n436) );
  CAOR2X1 U507 ( .A(\reg_mem[29][10] ), .B(n2418), .C(n2421), .D(n180), .Z(
        n437) );
  CAOR2X1 U508 ( .A(\reg_mem[29][9] ), .B(n2418), .C(n2422), .D(n181), .Z(n438) );
  CAOR2X1 U509 ( .A(\reg_mem[29][8] ), .B(n2418), .C(n2424), .D(n182), .Z(n439) );
  CAOR2X1 U510 ( .A(\reg_mem[29][7] ), .B(n2418), .C(n2422), .D(n183), .Z(n440) );
  CAOR2X1 U511 ( .A(\reg_mem[29][6] ), .B(n2418), .C(n2421), .D(n184), .Z(n441) );
  CAOR2X1 U512 ( .A(\reg_mem[29][5] ), .B(n2418), .C(n2422), .D(n185), .Z(n442) );
  CAOR2X1 U513 ( .A(\reg_mem[29][4] ), .B(n2418), .C(n2422), .D(n186), .Z(n443) );
  CAOR2X1 U514 ( .A(\reg_mem[29][3] ), .B(n2418), .C(n2421), .D(n187), .Z(n444) );
  CAOR2X1 U515 ( .A(\reg_mem[29][2] ), .B(n2418), .C(n2421), .D(n188), .Z(n445) );
  CAOR2X1 U516 ( .A(\reg_mem[29][1] ), .B(n2418), .C(n2423), .D(n189), .Z(n446) );
  CAOR2X1 U517 ( .A(\reg_mem[29][0] ), .B(n2418), .C(n2422), .D(n190), .Z(n447) );
  CAOR2X1 U518 ( .A(\reg_mem[28][31] ), .B(n2409), .C(n2417), .D(n2269), .Z(
        n448) );
  CAOR2X1 U519 ( .A(\reg_mem[28][30] ), .B(n2409), .C(n2416), .D(n2267), .Z(
        n449) );
  CAOR2X1 U520 ( .A(\reg_mem[28][29] ), .B(n2409), .C(n2417), .D(n2265), .Z(
        n450) );
  CAOR2X1 U521 ( .A(\reg_mem[28][28] ), .B(n2409), .C(n2417), .D(n2263), .Z(
        n451) );
  CAOR2X1 U522 ( .A(\reg_mem[28][27] ), .B(n2409), .C(n2416), .D(n2261), .Z(
        n452) );
  CAOR2X1 U523 ( .A(\reg_mem[28][26] ), .B(n2409), .C(n2416), .D(n2259), .Z(
        n453) );
  CAOR2X1 U524 ( .A(\reg_mem[28][25] ), .B(n2409), .C(n2415), .D(n2257), .Z(
        n454) );
  CAOR2X1 U525 ( .A(\reg_mem[28][24] ), .B(n2409), .C(n2415), .D(n2255), .Z(
        n455) );
  CAOR2X1 U526 ( .A(\reg_mem[28][23] ), .B(n197), .C(n2414), .D(n2253), .Z(
        n456) );
  CAOR2X1 U527 ( .A(\reg_mem[28][22] ), .B(n197), .C(n2413), .D(n2251), .Z(
        n457) );
  CAOR2X1 U528 ( .A(\reg_mem[28][21] ), .B(n1515), .C(n2415), .D(n2249), .Z(
        n458) );
  CAOR2X1 U529 ( .A(\reg_mem[28][20] ), .B(n1515), .C(n2415), .D(n2247), .Z(
        n459) );
  CAOR2X1 U530 ( .A(\reg_mem[28][19] ), .B(n1515), .C(n2414), .D(n2245), .Z(
        n460) );
  CAOR2X1 U531 ( .A(\reg_mem[28][18] ), .B(n1515), .C(n2413), .D(n2243), .Z(
        n461) );
  CAOR2X1 U532 ( .A(\reg_mem[28][17] ), .B(n1515), .C(n2414), .D(n2241), .Z(
        n462) );
  CAOR2X1 U533 ( .A(\reg_mem[28][16] ), .B(n1515), .C(n2414), .D(n2239), .Z(
        n463) );
  CAOR2X1 U534 ( .A(\reg_mem[28][15] ), .B(n1515), .C(n2413), .D(n2237), .Z(
        n464) );
  CAOR2X1 U535 ( .A(\reg_mem[28][14] ), .B(n1515), .C(n2413), .D(n2235), .Z(
        n465) );
  CAOR2X1 U536 ( .A(\reg_mem[28][13] ), .B(n1515), .C(n2412), .D(net83055), 
        .Z(n466) );
  CAOR2X1 U537 ( .A(\reg_mem[28][12] ), .B(n1515), .C(n2411), .D(n2233), .Z(
        n467) );
  CAOR2X1 U538 ( .A(\reg_mem[28][11] ), .B(n1515), .C(n2412), .D(net83059), 
        .Z(n468) );
  CAOR2X1 U539 ( .A(\reg_mem[28][10] ), .B(n1515), .C(n2412), .D(n2231), .Z(
        n469) );
  CAOR2X1 U540 ( .A(\reg_mem[28][9] ), .B(n1515), .C(n2411), .D(n2229), .Z(
        n470) );
  CAOR2X1 U541 ( .A(\reg_mem[28][8] ), .B(n1515), .C(n2411), .D(n2227), .Z(
        n471) );
  CAOR2X1 U542 ( .A(\reg_mem[28][7] ), .B(n1515), .C(n2410), .D(n2225), .Z(
        n472) );
  CAOR2X1 U543 ( .A(\reg_mem[28][6] ), .B(n1515), .C(n1514), .D(n2223), .Z(
        n473) );
  CAOR2X1 U544 ( .A(\reg_mem[28][5] ), .B(n1515), .C(n2410), .D(n2221), .Z(
        n474) );
  CAOR2X1 U545 ( .A(\reg_mem[28][4] ), .B(n1515), .C(n2410), .D(net83073), .Z(
        n475) );
  CAOR2X1 U546 ( .A(\reg_mem[28][3] ), .B(n1515), .C(n1514), .D(n2219), .Z(
        n476) );
  CAOR2X1 U547 ( .A(\reg_mem[28][2] ), .B(n1515), .C(n1514), .D(net83077), .Z(
        n477) );
  CAOR2X1 U548 ( .A(\reg_mem[28][1] ), .B(n1515), .C(n2417), .D(n2217), .Z(
        n478) );
  CAOR2X1 U549 ( .A(\reg_mem[28][0] ), .B(n1515), .C(n2416), .D(n2215), .Z(
        n479) );
  CAOR2X1 U550 ( .A(\reg_mem[27][31] ), .B(n2403), .C(n2405), .D(n2268), .Z(
        n480) );
  CAOR2X1 U551 ( .A(\reg_mem[27][30] ), .B(n2403), .C(n2405), .D(n2266), .Z(
        n481) );
  CAOR2X1 U552 ( .A(\reg_mem[27][29] ), .B(n2403), .C(n2408), .D(n2264), .Z(
        n482) );
  CAOR2X1 U553 ( .A(\reg_mem[27][28] ), .B(n2403), .C(n2408), .D(n2262), .Z(
        n483) );
  CAOR2X1 U554 ( .A(\reg_mem[27][27] ), .B(n2403), .C(n2408), .D(n2260), .Z(
        n484) );
  CAOR2X1 U555 ( .A(\reg_mem[27][26] ), .B(n2403), .C(n2406), .D(n2258), .Z(
        n485) );
  CAOR2X1 U556 ( .A(\reg_mem[27][25] ), .B(n2403), .C(n2408), .D(n2256), .Z(
        n486) );
  CAOR2X1 U557 ( .A(\reg_mem[27][24] ), .B(n2403), .C(n2408), .D(n2254), .Z(
        n487) );
  CAOR2X1 U558 ( .A(\reg_mem[27][23] ), .B(n199), .C(n2407), .D(n2252), .Z(
        n488) );
  CAOR2X1 U559 ( .A(\reg_mem[27][22] ), .B(n199), .C(n2407), .D(n2250), .Z(
        n489) );
  CAOR2X1 U560 ( .A(\reg_mem[27][21] ), .B(n1503), .C(n2408), .D(n2248), .Z(
        n490) );
  CAOR2X1 U561 ( .A(\reg_mem[27][20] ), .B(n1503), .C(n2408), .D(n2246), .Z(
        n491) );
  CAOR2X1 U562 ( .A(\reg_mem[27][19] ), .B(n1503), .C(n2406), .D(n2244), .Z(
        n492) );
  CAOR2X1 U563 ( .A(\reg_mem[27][18] ), .B(n1503), .C(n2407), .D(n2242), .Z(
        n493) );
  CAOR2X1 U564 ( .A(\reg_mem[27][17] ), .B(n1503), .C(n2405), .D(n2240), .Z(
        n494) );
  CAOR2X1 U565 ( .A(\reg_mem[27][16] ), .B(n1503), .C(n2407), .D(n2238), .Z(
        n495) );
  CAOR2X1 U566 ( .A(\reg_mem[27][15] ), .B(n1503), .C(n2407), .D(n2236), .Z(
        n496) );
  CAOR2X1 U567 ( .A(\reg_mem[27][14] ), .B(n1503), .C(n2407), .D(n2234), .Z(
        n497) );
  CAOR2X1 U568 ( .A(\reg_mem[27][13] ), .B(n1503), .C(n2406), .D(net83054), 
        .Z(n498) );
  CAOR2X1 U569 ( .A(\reg_mem[27][12] ), .B(n1503), .C(n2405), .D(n2232), .Z(
        n499) );
  CAOR2X1 U570 ( .A(\reg_mem[27][11] ), .B(n1503), .C(n2406), .D(net83058), 
        .Z(n500) );
  CAOR2X1 U571 ( .A(\reg_mem[27][10] ), .B(n1503), .C(n2406), .D(n2230), .Z(
        n501) );
  CAOR2X1 U572 ( .A(\reg_mem[27][9] ), .B(n1503), .C(n2405), .D(n2228), .Z(
        n502) );
  CAOR2X1 U573 ( .A(\reg_mem[27][8] ), .B(n1503), .C(n2405), .D(n2226), .Z(
        n503) );
  CAOR2X1 U574 ( .A(\reg_mem[27][7] ), .B(n1503), .C(n2404), .D(n2224), .Z(
        n504) );
  CAOR2X1 U575 ( .A(\reg_mem[27][6] ), .B(n1503), .C(n1502), .D(n2222), .Z(
        n505) );
  CAOR2X1 U576 ( .A(\reg_mem[27][5] ), .B(n1503), .C(n2404), .D(n2220), .Z(
        n506) );
  CAOR2X1 U577 ( .A(\reg_mem[27][4] ), .B(n1503), .C(n2404), .D(net83072), .Z(
        n507) );
  CAOR2X1 U578 ( .A(\reg_mem[27][3] ), .B(n1503), .C(n1502), .D(n2218), .Z(
        n508) );
  CAOR2X1 U579 ( .A(\reg_mem[27][2] ), .B(n1503), .C(n1502), .D(net83076), .Z(
        n509) );
  CAOR2X1 U580 ( .A(\reg_mem[27][1] ), .B(n1503), .C(n2406), .D(n2216), .Z(
        n510) );
  CAOR2X1 U581 ( .A(\reg_mem[27][0] ), .B(n1503), .C(n2406), .D(n2214), .Z(
        n511) );
  CAOR2X1 U582 ( .A(\reg_mem[26][31] ), .B(n1501), .C(n2402), .D(n159), .Z(
        n512) );
  CAOR2X1 U583 ( .A(\reg_mem[26][30] ), .B(n1501), .C(n2401), .D(n160), .Z(
        n513) );
  CAOR2X1 U584 ( .A(\reg_mem[26][29] ), .B(n1501), .C(n2402), .D(n161), .Z(
        n514) );
  CAOR2X1 U585 ( .A(\reg_mem[26][28] ), .B(n1501), .C(n2401), .D(n162), .Z(
        n515) );
  CAOR2X1 U586 ( .A(\reg_mem[26][27] ), .B(n1501), .C(n2401), .D(n163), .Z(
        n516) );
  CAOR2X1 U588 ( .A(\reg_mem[26][25] ), .B(n1501), .C(n1500), .D(n165), .Z(
        n518) );
  CAOR2X1 U589 ( .A(\reg_mem[26][24] ), .B(n1501), .C(n1500), .D(n166), .Z(
        n519) );
  CAOR2X1 U590 ( .A(\reg_mem[26][23] ), .B(n2398), .C(n1500), .D(n167), .Z(
        n520) );
  CAOR2X1 U591 ( .A(\reg_mem[26][22] ), .B(n2398), .C(n1500), .D(n168), .Z(
        n521) );
  CAOR2X1 U592 ( .A(\reg_mem[26][21] ), .B(n2398), .C(n2402), .D(n169), .Z(
        n522) );
  CAOR2X1 U593 ( .A(\reg_mem[26][20] ), .B(n2398), .C(n2401), .D(n170), .Z(
        n523) );
  CAOR2X1 U594 ( .A(\reg_mem[26][19] ), .B(n2398), .C(n2402), .D(n171), .Z(
        n524) );
  CAOR2X1 U595 ( .A(\reg_mem[26][18] ), .B(n2398), .C(n2401), .D(n172), .Z(
        n525) );
  CAOR2X1 U596 ( .A(\reg_mem[26][17] ), .B(n2398), .C(n2402), .D(n173), .Z(
        n526) );
  CAOR2X1 U597 ( .A(\reg_mem[26][16] ), .B(n2398), .C(n2402), .D(n174), .Z(
        n527) );
  CAOR2X1 U598 ( .A(\reg_mem[26][15] ), .B(n2398), .C(n2401), .D(n175), .Z(
        n528) );
  CAOR2X1 U599 ( .A(\reg_mem[26][14] ), .B(n2398), .C(n2401), .D(n176), .Z(
        n529) );
  CAOR2X1 U600 ( .A(\reg_mem[26][13] ), .B(n2398), .C(n2400), .D(n177), .Z(
        n530) );
  CAOR2X1 U601 ( .A(\reg_mem[26][12] ), .B(n2398), .C(n2399), .D(n178), .Z(
        n531) );
  CAOR2X1 U602 ( .A(\reg_mem[26][11] ), .B(n2397), .C(n2400), .D(n179), .Z(
        n532) );
  CAOR2X1 U603 ( .A(\reg_mem[26][10] ), .B(n2397), .C(n2399), .D(n180), .Z(
        n533) );
  CAOR2X1 U604 ( .A(\reg_mem[26][9] ), .B(n2397), .C(n2400), .D(n181), .Z(n534) );
  CAOR2X1 U605 ( .A(\reg_mem[26][8] ), .B(n2397), .C(n2399), .D(n182), .Z(n535) );
  CAOR2X1 U606 ( .A(\reg_mem[26][7] ), .B(n2397), .C(n2400), .D(n183), .Z(n536) );
  CAOR2X1 U607 ( .A(\reg_mem[26][6] ), .B(n2397), .C(n2399), .D(n184), .Z(n537) );
  CAOR2X1 U608 ( .A(\reg_mem[26][5] ), .B(n2397), .C(n2400), .D(n185), .Z(n538) );
  CAOR2X1 U609 ( .A(\reg_mem[26][4] ), .B(n2397), .C(n2400), .D(n186), .Z(n539) );
  CAOR2X1 U610 ( .A(\reg_mem[26][3] ), .B(n2397), .C(n2399), .D(n187), .Z(n540) );
  CAOR2X1 U611 ( .A(\reg_mem[26][2] ), .B(n2397), .C(n2399), .D(n188), .Z(n541) );
  CAOR2X1 U612 ( .A(\reg_mem[26][1] ), .B(n2397), .C(n2402), .D(n189), .Z(n542) );
  CAOR2X1 U613 ( .A(\reg_mem[26][0] ), .B(n2397), .C(n1500), .D(n190), .Z(n543) );
  CAOR2X1 U614 ( .A(\reg_mem[25][31] ), .B(n2388), .C(n2396), .D(n2269), .Z(
        n544) );
  CAOR2X1 U615 ( .A(\reg_mem[25][30] ), .B(n2388), .C(n2395), .D(n2267), .Z(
        n545) );
  CAOR2X1 U616 ( .A(\reg_mem[25][29] ), .B(n2388), .C(n2396), .D(n2265), .Z(
        n546) );
  CAOR2X1 U617 ( .A(\reg_mem[25][28] ), .B(n2388), .C(n2396), .D(n2263), .Z(
        n547) );
  CAOR2X1 U618 ( .A(\reg_mem[25][27] ), .B(n2388), .C(n2395), .D(n2261), .Z(
        n548) );
  CAOR2X1 U619 ( .A(\reg_mem[25][26] ), .B(n2388), .C(n2395), .D(n2259), .Z(
        n549) );
  CAOR2X1 U620 ( .A(\reg_mem[25][25] ), .B(n2388), .C(n2394), .D(n2257), .Z(
        n550) );
  CAOR2X1 U621 ( .A(\reg_mem[25][24] ), .B(n2388), .C(n2394), .D(n2255), .Z(
        n551) );
  CAOR2X1 U622 ( .A(\reg_mem[25][23] ), .B(n1513), .C(n2393), .D(n2253), .Z(
        n552) );
  CAOR2X1 U623 ( .A(\reg_mem[25][22] ), .B(n1513), .C(n2392), .D(n2251), .Z(
        n553) );
  CAOR2X1 U624 ( .A(\reg_mem[25][21] ), .B(n1513), .C(n2394), .D(n2249), .Z(
        n554) );
  CAOR2X1 U625 ( .A(\reg_mem[25][20] ), .B(n1513), .C(n2394), .D(n2247), .Z(
        n555) );
  CAOR2X1 U626 ( .A(\reg_mem[25][19] ), .B(n1513), .C(n2393), .D(n2245), .Z(
        n556) );
  CAOR2X1 U627 ( .A(\reg_mem[25][18] ), .B(n1513), .C(n2392), .D(n2243), .Z(
        n557) );
  CAOR2X1 U628 ( .A(\reg_mem[25][17] ), .B(n1513), .C(n2393), .D(n2241), .Z(
        n558) );
  CAOR2X1 U629 ( .A(\reg_mem[25][16] ), .B(n1513), .C(n2393), .D(n2239), .Z(
        n559) );
  CAOR2X1 U630 ( .A(\reg_mem[25][15] ), .B(n1513), .C(n2392), .D(n2237), .Z(
        n560) );
  CAOR2X1 U631 ( .A(\reg_mem[25][14] ), .B(n1513), .C(n2392), .D(n2235), .Z(
        n561) );
  CAOR2X1 U632 ( .A(\reg_mem[25][13] ), .B(n1513), .C(n2391), .D(net83055), 
        .Z(n562) );
  CAOR2X1 U633 ( .A(\reg_mem[25][12] ), .B(n1513), .C(n1512), .D(n2233), .Z(
        n563) );
  CAOR2X1 U634 ( .A(\reg_mem[25][11] ), .B(n1513), .C(n2391), .D(net83059), 
        .Z(n564) );
  CAOR2X1 U635 ( .A(\reg_mem[25][10] ), .B(n1513), .C(n2391), .D(n2231), .Z(
        n565) );
  CAOR2X1 U636 ( .A(\reg_mem[25][9] ), .B(n1513), .C(n1512), .D(n2229), .Z(
        n566) );
  CAOR2X1 U637 ( .A(\reg_mem[25][8] ), .B(n1513), .C(n1512), .D(n2227), .Z(
        n567) );
  CAOR2X1 U638 ( .A(\reg_mem[25][7] ), .B(n1513), .C(n2390), .D(n2225), .Z(
        n568) );
  CAOR2X1 U639 ( .A(\reg_mem[25][6] ), .B(n1513), .C(n2389), .D(n2223), .Z(
        n569) );
  CAOR2X1 U640 ( .A(\reg_mem[25][5] ), .B(n1513), .C(n2390), .D(n2221), .Z(
        n570) );
  CAOR2X1 U641 ( .A(\reg_mem[25][4] ), .B(n1513), .C(n2390), .D(net83073), .Z(
        n571) );
  CAOR2X1 U642 ( .A(\reg_mem[25][3] ), .B(n1513), .C(n2389), .D(n2219), .Z(
        n572) );
  CAOR2X1 U643 ( .A(\reg_mem[25][2] ), .B(n1513), .C(n2389), .D(net83077), .Z(
        n573) );
  CAOR2X1 U644 ( .A(\reg_mem[25][1] ), .B(n1513), .C(n2396), .D(n2217), .Z(
        n574) );
  CAOR2X1 U645 ( .A(\reg_mem[25][0] ), .B(n1513), .C(n2395), .D(n2215), .Z(
        n575) );
  CAOR2X1 U646 ( .A(\reg_mem[24][31] ), .B(n2379), .C(n2387), .D(n2268), .Z(
        n576) );
  CAOR2X1 U647 ( .A(\reg_mem[24][30] ), .B(n2379), .C(n2386), .D(n2266), .Z(
        n577) );
  CAOR2X1 U648 ( .A(\reg_mem[24][29] ), .B(n2379), .C(n2387), .D(n2264), .Z(
        n578) );
  CAOR2X1 U649 ( .A(\reg_mem[24][28] ), .B(n2379), .C(n2387), .D(n2262), .Z(
        n579) );
  CAOR2X1 U650 ( .A(\reg_mem[24][27] ), .B(n2379), .C(n2386), .D(n2260), .Z(
        n580) );
  CAOR2X1 U651 ( .A(\reg_mem[24][26] ), .B(n2379), .C(n2386), .D(n2258), .Z(
        n581) );
  CAOR2X1 U652 ( .A(\reg_mem[24][25] ), .B(n2379), .C(n2385), .D(n2256), .Z(
        n582) );
  CAOR2X1 U653 ( .A(\reg_mem[24][24] ), .B(n2379), .C(n2385), .D(n2254), .Z(
        n583) );
  CAOR2X1 U654 ( .A(\reg_mem[24][23] ), .B(n1511), .C(n2384), .D(n2252), .Z(
        n584) );
  CAOR2X1 U655 ( .A(\reg_mem[24][22] ), .B(n1511), .C(n2383), .D(n2250), .Z(
        n585) );
  CAOR2X1 U656 ( .A(\reg_mem[24][21] ), .B(n1511), .C(n2385), .D(n2248), .Z(
        n586) );
  CAOR2X1 U657 ( .A(\reg_mem[24][20] ), .B(n1511), .C(n2385), .D(n2246), .Z(
        n587) );
  CAOR2X1 U658 ( .A(\reg_mem[24][19] ), .B(n1511), .C(n2384), .D(n2244), .Z(
        n588) );
  CAOR2X1 U659 ( .A(\reg_mem[24][18] ), .B(n1511), .C(n2383), .D(n2242), .Z(
        n589) );
  CAOR2X1 U660 ( .A(\reg_mem[24][17] ), .B(n1511), .C(n2384), .D(n2240), .Z(
        n590) );
  CAOR2X1 U661 ( .A(\reg_mem[24][16] ), .B(n1511), .C(n2384), .D(n2238), .Z(
        n591) );
  CAOR2X1 U662 ( .A(\reg_mem[24][15] ), .B(n1511), .C(n2383), .D(n2236), .Z(
        n592) );
  CAOR2X1 U663 ( .A(\reg_mem[24][14] ), .B(n1511), .C(n2383), .D(n2234), .Z(
        n593) );
  CAOR2X1 U664 ( .A(\reg_mem[24][13] ), .B(n1511), .C(n2382), .D(net83054), 
        .Z(n594) );
  CAOR2X1 U665 ( .A(\reg_mem[24][12] ), .B(n1511), .C(n1510), .D(n2232), .Z(
        n595) );
  CAOR2X1 U666 ( .A(\reg_mem[24][11] ), .B(n1511), .C(n2382), .D(net83058), 
        .Z(n596) );
  CAOR2X1 U667 ( .A(\reg_mem[24][10] ), .B(n1511), .C(n2382), .D(n2230), .Z(
        n597) );
  CAOR2X1 U668 ( .A(\reg_mem[24][9] ), .B(n1511), .C(n1510), .D(n2228), .Z(
        n598) );
  CAOR2X1 U669 ( .A(\reg_mem[24][8] ), .B(n1511), .C(n1510), .D(n2226), .Z(
        n599) );
  CAOR2X1 U670 ( .A(\reg_mem[24][7] ), .B(n1511), .C(n2381), .D(n2224), .Z(
        n600) );
  CAOR2X1 U671 ( .A(\reg_mem[24][6] ), .B(n1511), .C(n2380), .D(n2222), .Z(
        n601) );
  CAOR2X1 U672 ( .A(\reg_mem[24][5] ), .B(n1511), .C(n2381), .D(n2220), .Z(
        n602) );
  CAOR2X1 U673 ( .A(\reg_mem[24][4] ), .B(n1511), .C(n2381), .D(net83072), .Z(
        n603) );
  CAOR2X1 U674 ( .A(\reg_mem[24][3] ), .B(n1511), .C(n2380), .D(n2218), .Z(
        n604) );
  CAOR2X1 U675 ( .A(\reg_mem[24][2] ), .B(n1511), .C(n2380), .D(net83076), .Z(
        n605) );
  CAOR2X1 U676 ( .A(\reg_mem[24][1] ), .B(n1511), .C(n2387), .D(n2216), .Z(
        n606) );
  CAOR2X1 U677 ( .A(\reg_mem[24][0] ), .B(n1511), .C(n2386), .D(n2214), .Z(
        n607) );
  CAOR2X1 U678 ( .A(\reg_mem[23][31] ), .B(n2374), .C(n2377), .D(n159), .Z(
        n608) );
  CAOR2X1 U679 ( .A(\reg_mem[23][30] ), .B(n2374), .C(n2375), .D(n160), .Z(
        n609) );
  CAOR2X1 U680 ( .A(\reg_mem[23][29] ), .B(n2374), .C(n2377), .D(n161), .Z(
        n610) );
  CAOR2X1 U681 ( .A(\reg_mem[23][28] ), .B(n2374), .C(n2376), .D(n162), .Z(
        n611) );
  CAOR2X1 U682 ( .A(\reg_mem[23][27] ), .B(n2374), .C(n2376), .D(n163), .Z(
        n612) );
  CAOR2X1 U683 ( .A(\reg_mem[23][26] ), .B(n2374), .C(n2377), .D(n164), .Z(
        n613) );
  CAOR2X1 U684 ( .A(\reg_mem[23][25] ), .B(n2374), .C(n2375), .D(n165), .Z(
        n614) );
  CAOR2X1 U685 ( .A(\reg_mem[23][24] ), .B(n2374), .C(n2376), .D(n166), .Z(
        n615) );
  CAOR2X1 U686 ( .A(\reg_mem[23][23] ), .B(n2373), .C(n2376), .D(n167), .Z(
        n616) );
  CAOR2X1 U687 ( .A(\reg_mem[23][22] ), .B(n2373), .C(n2377), .D(n168), .Z(
        n617) );
  CAOR2X1 U688 ( .A(\reg_mem[23][21] ), .B(n2373), .C(n2377), .D(n169), .Z(
        n618) );
  CAOR2X1 U689 ( .A(\reg_mem[23][20] ), .B(n2373), .C(n2375), .D(n170), .Z(
        n619) );
  CAOR2X1 U690 ( .A(\reg_mem[23][19] ), .B(n2373), .C(n2377), .D(n171), .Z(
        n620) );
  CAOR2X1 U691 ( .A(\reg_mem[23][18] ), .B(n2373), .C(n2375), .D(n172), .Z(
        n621) );
  CAOR2X1 U692 ( .A(\reg_mem[23][17] ), .B(n2373), .C(n2376), .D(n173), .Z(
        n622) );
  CAOR2X1 U693 ( .A(\reg_mem[23][16] ), .B(n2373), .C(n2375), .D(n174), .Z(
        n623) );
  CAOR2X1 U694 ( .A(\reg_mem[23][15] ), .B(n2373), .C(n2377), .D(n175), .Z(
        n624) );
  CAOR2X1 U695 ( .A(\reg_mem[23][14] ), .B(n2373), .C(n2377), .D(n176), .Z(
        n625) );
  CAOR2X1 U696 ( .A(\reg_mem[23][13] ), .B(n2373), .C(n2376), .D(n177), .Z(
        n626) );
  CAOR2X1 U697 ( .A(\reg_mem[23][12] ), .B(n2373), .C(n2375), .D(n178), .Z(
        n627) );
  CAOR2X1 U698 ( .A(\reg_mem[23][11] ), .B(n2372), .C(n2377), .D(n179), .Z(
        n628) );
  CAOR2X1 U699 ( .A(\reg_mem[23][10] ), .B(n2372), .C(n2377), .D(n180), .Z(
        n629) );
  CAOR2X1 U700 ( .A(\reg_mem[23][9] ), .B(n2372), .C(n2375), .D(n181), .Z(n630) );
  CAOR2X1 U701 ( .A(\reg_mem[23][8] ), .B(n2372), .C(n2376), .D(n182), .Z(n631) );
  CAOR2X1 U702 ( .A(\reg_mem[23][7] ), .B(n2372), .C(n2376), .D(n183), .Z(n632) );
  CAOR2X1 U703 ( .A(\reg_mem[23][6] ), .B(n2372), .C(n2375), .D(n184), .Z(n633) );
  CAOR2X1 U704 ( .A(\reg_mem[23][5] ), .B(n2372), .C(n2376), .D(n185), .Z(n634) );
  CAOR2X1 U705 ( .A(\reg_mem[23][4] ), .B(n2372), .C(n2376), .D(n186), .Z(n635) );
  CAOR2X1 U706 ( .A(\reg_mem[23][3] ), .B(n2372), .C(n2375), .D(n187), .Z(n636) );
  CAOR2X1 U707 ( .A(\reg_mem[23][2] ), .B(n2372), .C(n2375), .D(n188), .Z(n637) );
  CAOR2X1 U708 ( .A(\reg_mem[23][1] ), .B(n2372), .C(n2375), .D(n189), .Z(n638) );
  CAOR2X1 U709 ( .A(\reg_mem[23][0] ), .B(n2372), .C(n2377), .D(n190), .Z(n639) );
  CAOR2X1 U710 ( .A(\reg_mem[22][31] ), .B(n2363), .C(n2370), .D(n2269), .Z(
        n640) );
  CAOR2X1 U711 ( .A(\reg_mem[22][30] ), .B(n2363), .C(n2366), .D(n2267), .Z(
        n641) );
  CAOR2X1 U712 ( .A(\reg_mem[22][29] ), .B(n2363), .C(n2369), .D(n2265), .Z(
        n642) );
  CAOR2X1 U713 ( .A(\reg_mem[22][28] ), .B(n2363), .C(n2368), .D(n2263), .Z(
        n643) );
  CAOR2X1 U714 ( .A(\reg_mem[22][27] ), .B(n2363), .C(n2365), .D(n2261), .Z(
        n644) );
  CAOR2X1 U715 ( .A(\reg_mem[22][26] ), .B(n2363), .C(n2364), .D(n2259), .Z(
        n645) );
  CAOR2X1 U716 ( .A(\reg_mem[22][25] ), .B(n1529), .C(n2371), .D(n2257), .Z(
        n646) );
  CAOR2X1 U717 ( .A(\reg_mem[22][24] ), .B(n2363), .C(n2370), .D(n2255), .Z(
        n647) );
  CAOR2X1 U718 ( .A(\reg_mem[22][23] ), .B(n1529), .C(n2371), .D(n2253), .Z(
        n648) );
  CAOR2X1 U719 ( .A(\reg_mem[22][22] ), .B(n1529), .C(n2371), .D(n2251), .Z(
        n649) );
  CAOR2X1 U720 ( .A(\reg_mem[22][21] ), .B(n1529), .C(n2370), .D(n2249), .Z(
        n650) );
  CAOR2X1 U721 ( .A(\reg_mem[22][20] ), .B(n1529), .C(n2370), .D(n2247), .Z(
        n651) );
  CAOR2X1 U722 ( .A(\reg_mem[22][19] ), .B(n1529), .C(n2369), .D(n2245), .Z(
        n652) );
  CAOR2X1 U723 ( .A(\reg_mem[22][18] ), .B(n1529), .C(n2368), .D(n2243), .Z(
        n653) );
  CAOR2X1 U724 ( .A(\reg_mem[22][17] ), .B(n1529), .C(n2369), .D(n2241), .Z(
        n654) );
  CAOR2X1 U725 ( .A(\reg_mem[22][16] ), .B(n1529), .C(n2369), .D(n2239), .Z(
        n655) );
  CAOR2X1 U726 ( .A(\reg_mem[22][15] ), .B(n1529), .C(n2368), .D(n2237), .Z(
        n656) );
  CAOR2X1 U727 ( .A(\reg_mem[22][14] ), .B(n1529), .C(n2368), .D(n2235), .Z(
        n657) );
  CAOR2X1 U728 ( .A(\reg_mem[22][13] ), .B(n1529), .C(n2367), .D(net83055), 
        .Z(n658) );
  CAOR2X1 U729 ( .A(\reg_mem[22][12] ), .B(n1529), .C(n2366), .D(n2233), .Z(
        n659) );
  CAOR2X1 U730 ( .A(\reg_mem[22][11] ), .B(n2363), .C(n2367), .D(net83059), 
        .Z(n660) );
  CAOR2X1 U731 ( .A(\reg_mem[22][10] ), .B(n2363), .C(n2367), .D(n2231), .Z(
        n661) );
  CAOR2X1 U732 ( .A(\reg_mem[22][9] ), .B(n2363), .C(n2366), .D(n2229), .Z(
        n662) );
  CAOR2X1 U733 ( .A(\reg_mem[22][8] ), .B(n2363), .C(n2366), .D(n2227), .Z(
        n663) );
  CAOR2X1 U734 ( .A(\reg_mem[22][7] ), .B(n2363), .C(n2365), .D(n2225), .Z(
        n664) );
  CAOR2X1 U735 ( .A(\reg_mem[22][6] ), .B(n2363), .C(n2364), .D(n2223), .Z(
        n665) );
  CAOR2X1 U736 ( .A(\reg_mem[22][5] ), .B(n2363), .C(n2365), .D(n2221), .Z(
        n666) );
  CAOR2X1 U737 ( .A(\reg_mem[22][4] ), .B(n2363), .C(n2365), .D(net83073), .Z(
        n667) );
  CAOR2X1 U738 ( .A(\reg_mem[22][3] ), .B(n2363), .C(n2364), .D(n2219), .Z(
        n668) );
  CAOR2X1 U739 ( .A(\reg_mem[22][2] ), .B(n2363), .C(n2364), .D(net83077), .Z(
        n669) );
  CAOR2X1 U740 ( .A(\reg_mem[22][1] ), .B(n2363), .C(n2371), .D(n2217), .Z(
        n670) );
  CAOR2X1 U741 ( .A(\reg_mem[22][0] ), .B(n2363), .C(n2367), .D(n2215), .Z(
        n671) );
  CAOR2X1 U742 ( .A(\reg_mem[21][31] ), .B(n2357), .C(n2362), .D(n2268), .Z(
        n672) );
  CAOR2X1 U743 ( .A(\reg_mem[21][30] ), .B(n2357), .C(n2360), .D(n2266), .Z(
        n673) );
  CAOR2X1 U744 ( .A(\reg_mem[21][29] ), .B(n2357), .C(n2361), .D(n2264), .Z(
        n674) );
  CAOR2X1 U745 ( .A(\reg_mem[21][28] ), .B(n2357), .C(n2360), .D(n2262), .Z(
        n675) );
  CAOR2X1 U746 ( .A(\reg_mem[21][27] ), .B(n2357), .C(n2362), .D(n2260), .Z(
        n676) );
  CAOR2X1 U747 ( .A(\reg_mem[21][26] ), .B(n2357), .C(n2361), .D(n2258), .Z(
        n677) );
  CAOR2X1 U748 ( .A(\reg_mem[21][25] ), .B(n2357), .C(n2362), .D(n2256), .Z(
        n678) );
  CAOR2X1 U749 ( .A(\reg_mem[21][24] ), .B(n2357), .C(n2362), .D(n2254), .Z(
        n679) );
  CAOR2X1 U750 ( .A(\reg_mem[21][23] ), .B(n1521), .C(n2361), .D(n2252), .Z(
        n680) );
  CAOR2X1 U751 ( .A(\reg_mem[21][22] ), .B(n1521), .C(n2360), .D(n2250), .Z(
        n681) );
  CAOR2X1 U752 ( .A(\reg_mem[21][21] ), .B(n1521), .C(n2362), .D(n2248), .Z(
        n682) );
  CAOR2X1 U753 ( .A(\reg_mem[21][20] ), .B(n1521), .C(n2362), .D(n2246), .Z(
        n683) );
  CAOR2X1 U754 ( .A(\reg_mem[21][19] ), .B(n1521), .C(n2361), .D(n2244), .Z(
        n684) );
  CAOR2X1 U755 ( .A(\reg_mem[21][18] ), .B(n1521), .C(n2360), .D(n2242), .Z(
        n685) );
  CAOR2X1 U756 ( .A(\reg_mem[21][17] ), .B(n1521), .C(n2361), .D(n2240), .Z(
        n686) );
  CAOR2X1 U757 ( .A(\reg_mem[21][16] ), .B(n1521), .C(n2361), .D(n2238), .Z(
        n687) );
  CAOR2X1 U758 ( .A(\reg_mem[21][15] ), .B(n1521), .C(n2360), .D(n2236), .Z(
        n688) );
  CAOR2X1 U759 ( .A(\reg_mem[21][14] ), .B(n1521), .C(n2360), .D(n2234), .Z(
        n689) );
  CAOR2X1 U760 ( .A(\reg_mem[21][13] ), .B(n1521), .C(n2359), .D(net83054), 
        .Z(n690) );
  CAOR2X1 U761 ( .A(\reg_mem[21][12] ), .B(n1521), .C(n2358), .D(n2232), .Z(
        n691) );
  CAOR2X1 U762 ( .A(\reg_mem[21][11] ), .B(n1521), .C(n2359), .D(net83058), 
        .Z(n692) );
  CAOR2X1 U763 ( .A(\reg_mem[21][10] ), .B(n1521), .C(n2358), .D(n2230), .Z(
        n693) );
  CAOR2X1 U764 ( .A(\reg_mem[21][9] ), .B(n1521), .C(n2359), .D(n2228), .Z(
        n694) );
  CAOR2X1 U765 ( .A(\reg_mem[21][8] ), .B(n1521), .C(n2358), .D(n2226), .Z(
        n695) );
  CAOR2X1 U766 ( .A(\reg_mem[21][7] ), .B(n1521), .C(n2359), .D(n2224), .Z(
        n696) );
  CAOR2X1 U767 ( .A(\reg_mem[21][6] ), .B(n1521), .C(n2358), .D(n2222), .Z(
        n697) );
  CAOR2X1 U768 ( .A(\reg_mem[21][5] ), .B(n1521), .C(n2359), .D(n2220), .Z(
        n698) );
  CAOR2X1 U769 ( .A(\reg_mem[21][4] ), .B(n1521), .C(n2359), .D(net83072), .Z(
        n699) );
  CAOR2X1 U770 ( .A(\reg_mem[21][3] ), .B(n212), .C(n2358), .D(n2218), .Z(n700) );
  CAOR2X1 U771 ( .A(\reg_mem[21][2] ), .B(n212), .C(n2358), .D(net83076), .Z(
        n701) );
  CAOR2X1 U772 ( .A(\reg_mem[21][1] ), .B(n212), .C(n2362), .D(n2216), .Z(n702) );
  CAOR2X1 U773 ( .A(\reg_mem[21][0] ), .B(n212), .C(n2361), .D(n2214), .Z(n703) );
  CAOR2X1 U774 ( .A(\reg_mem[20][31] ), .B(n2351), .C(n2354), .D(n159), .Z(
        n704) );
  CAOR2X1 U775 ( .A(\reg_mem[20][30] ), .B(n2351), .C(n2356), .D(n160), .Z(
        n705) );
  CAOR2X1 U777 ( .A(\reg_mem[20][28] ), .B(n2351), .C(n2352), .D(n162), .Z(
        n707) );
  CAOR2X1 U778 ( .A(\reg_mem[20][27] ), .B(n2351), .C(n2356), .D(n163), .Z(
        n708) );
  CAOR2X1 U779 ( .A(\reg_mem[20][26] ), .B(n2351), .C(n2355), .D(n164), .Z(
        n709) );
  CAOR2X1 U780 ( .A(\reg_mem[20][25] ), .B(n2351), .C(n2356), .D(n165), .Z(
        n710) );
  CAOR2X1 U781 ( .A(\reg_mem[20][24] ), .B(n2351), .C(n2356), .D(n166), .Z(
        n711) );
  CAOR2X1 U782 ( .A(\reg_mem[20][23] ), .B(n1519), .C(n2355), .D(n167), .Z(
        n712) );
  CAOR2X1 U783 ( .A(\reg_mem[20][22] ), .B(n1519), .C(n2354), .D(n168), .Z(
        n713) );
  CAOR2X1 U784 ( .A(\reg_mem[20][21] ), .B(n1519), .C(n2356), .D(n169), .Z(
        n714) );
  CAOR2X1 U785 ( .A(\reg_mem[20][20] ), .B(n1519), .C(n2356), .D(n170), .Z(
        n715) );
  CAOR2X1 U786 ( .A(\reg_mem[20][19] ), .B(n1519), .C(n2355), .D(n171), .Z(
        n716) );
  CAOR2X1 U787 ( .A(\reg_mem[20][18] ), .B(n1519), .C(n2354), .D(n172), .Z(
        n717) );
  CAOR2X1 U788 ( .A(\reg_mem[20][17] ), .B(n1519), .C(n2355), .D(n173), .Z(
        n718) );
  CAOR2X1 U789 ( .A(\reg_mem[20][16] ), .B(n1519), .C(n2355), .D(n174), .Z(
        n719) );
  CAOR2X1 U790 ( .A(\reg_mem[20][15] ), .B(n1519), .C(n2354), .D(n175), .Z(
        n720) );
  CAOR2X1 U791 ( .A(\reg_mem[20][14] ), .B(n1519), .C(n2354), .D(n176), .Z(
        n721) );
  CAOR2X1 U792 ( .A(\reg_mem[20][13] ), .B(n1519), .C(n2353), .D(n177), .Z(
        n722) );
  CAOR2X1 U793 ( .A(\reg_mem[20][12] ), .B(n1519), .C(n2352), .D(n178), .Z(
        n723) );
  CAOR2X1 U794 ( .A(\reg_mem[20][11] ), .B(n1519), .C(n2353), .D(n179), .Z(
        n724) );
  CAOR2X1 U795 ( .A(\reg_mem[20][10] ), .B(n1519), .C(n2352), .D(n180), .Z(
        n725) );
  CAOR2X1 U796 ( .A(\reg_mem[20][9] ), .B(n1519), .C(n2354), .D(n181), .Z(n726) );
  CAOR2X1 U797 ( .A(\reg_mem[20][8] ), .B(n1519), .C(n2353), .D(n182), .Z(n727) );
  CAOR2X1 U798 ( .A(\reg_mem[20][7] ), .B(n1519), .C(n2353), .D(n183), .Z(n728) );
  CAOR2X1 U799 ( .A(\reg_mem[20][6] ), .B(n1519), .C(n2352), .D(n184), .Z(n729) );
  CAOR2X1 U800 ( .A(\reg_mem[20][5] ), .B(n1519), .C(n2353), .D(n185), .Z(n730) );
  CAOR2X1 U801 ( .A(\reg_mem[20][4] ), .B(n213), .C(n2353), .D(n186), .Z(n731)
         );
  CAOR2X1 U802 ( .A(\reg_mem[20][3] ), .B(n213), .C(n2352), .D(n187), .Z(n732)
         );
  CAOR2X1 U803 ( .A(\reg_mem[20][2] ), .B(n213), .C(n2352), .D(n188), .Z(n733)
         );
  CAOR2X1 U804 ( .A(\reg_mem[20][1] ), .B(n213), .C(n2356), .D(n189), .Z(n734)
         );
  CAOR2X1 U805 ( .A(\reg_mem[20][0] ), .B(n213), .C(n2355), .D(n190), .Z(n735)
         );
  CAOR2X1 U806 ( .A(\reg_mem[19][31] ), .B(net81901), .C(net81923), .D(n2269), 
        .Z(n736) );
  CAOR2X1 U807 ( .A(\reg_mem[19][30] ), .B(net81901), .C(net81917), .D(n2267), 
        .Z(n737) );
  CAOR2X1 U808 ( .A(\reg_mem[19][29] ), .B(net81901), .C(net81919), .D(n2265), 
        .Z(n738) );
  CAOR2X1 U809 ( .A(\reg_mem[19][28] ), .B(net81901), .C(net81917), .D(n2263), 
        .Z(n739) );
  CAOR2X1 U810 ( .A(\reg_mem[19][27] ), .B(net81901), .C(net81923), .D(n2261), 
        .Z(n740) );
  CAOR2X1 U811 ( .A(\reg_mem[19][26] ), .B(net81901), .C(net81919), .D(n2259), 
        .Z(n741) );
  CAOR2X1 U812 ( .A(\reg_mem[19][25] ), .B(net81901), .C(net81923), .D(n2257), 
        .Z(n742) );
  CAOR2X1 U813 ( .A(\reg_mem[19][24] ), .B(net81901), .C(net81923), .D(n2255), 
        .Z(n743) );
  CAOR2X1 U814 ( .A(\reg_mem[19][23] ), .B(n1517), .C(net81919), .D(n2253), 
        .Z(n744) );
  CAOR2X1 U815 ( .A(\reg_mem[19][22] ), .B(n1517), .C(net81917), .D(n2251), 
        .Z(n745) );
  CAOR2X1 U816 ( .A(\reg_mem[19][21] ), .B(n1517), .C(net81923), .D(n2249), 
        .Z(n746) );
  CAOR2X1 U817 ( .A(\reg_mem[19][20] ), .B(n1517), .C(net81923), .D(n2247), 
        .Z(n747) );
  CAOR2X1 U818 ( .A(\reg_mem[19][19] ), .B(n1517), .C(net81919), .D(n2245), 
        .Z(n748) );
  CAOR2X1 U819 ( .A(\reg_mem[19][18] ), .B(n1517), .C(net81917), .D(n2243), 
        .Z(n749) );
  CAOR2X1 U820 ( .A(\reg_mem[19][17] ), .B(n1517), .C(net81919), .D(n2241), 
        .Z(n750) );
  CAOR2X1 U821 ( .A(\reg_mem[19][16] ), .B(n1517), .C(net81919), .D(n2239), 
        .Z(n751) );
  CAOR2X1 U822 ( .A(\reg_mem[19][15] ), .B(n1517), .C(net81917), .D(n2237), 
        .Z(n752) );
  CAOR2X1 U823 ( .A(\reg_mem[19][14] ), .B(n1517), .C(net81917), .D(n2235), 
        .Z(n753) );
  CAOR2X1 U824 ( .A(\reg_mem[19][13] ), .B(n1517), .C(net81907), .D(net83055), 
        .Z(n754) );
  CAOR2X1 U825 ( .A(\reg_mem[19][12] ), .B(n1517), .C(net81905), .D(n2233), 
        .Z(n755) );
  CAOR2X1 U826 ( .A(\reg_mem[19][11] ), .B(n1517), .C(net81907), .D(net83059), 
        .Z(n756) );
  CAOR2X1 U827 ( .A(\reg_mem[19][10] ), .B(n1517), .C(net81905), .D(n2231), 
        .Z(n757) );
  CAOR2X1 U828 ( .A(\reg_mem[19][9] ), .B(n1517), .C(net81907), .D(n2229), .Z(
        n758) );
  CAOR2X1 U829 ( .A(\reg_mem[19][8] ), .B(n1517), .C(net81905), .D(n2227), .Z(
        n759) );
  CAOR2X1 U830 ( .A(\reg_mem[19][7] ), .B(n1517), .C(net81907), .D(n2225), .Z(
        n760) );
  CAOR2X1 U831 ( .A(\reg_mem[19][6] ), .B(n1517), .C(net81905), .D(n2223), .Z(
        n761) );
  CAOR2X1 U832 ( .A(\reg_mem[19][5] ), .B(n1517), .C(net81907), .D(n2221), .Z(
        n762) );
  CAOR2X1 U834 ( .A(\reg_mem[19][3] ), .B(n1517), .C(net81905), .D(n2219), .Z(
        n764) );
  CAOR2X1 U836 ( .A(\reg_mem[19][1] ), .B(n214), .C(net81923), .D(n2217), .Z(
        n766) );
  CAOR2X1 U837 ( .A(\reg_mem[19][0] ), .B(n214), .C(net81919), .D(n2215), .Z(
        n767) );
  CAOR2X1 U838 ( .A(\reg_mem[18][31] ), .B(net81941), .C(net81971), .D(n2268), 
        .Z(n768) );
  CAOR2X1 U839 ( .A(\reg_mem[18][30] ), .B(net81941), .C(n1506), .D(n2266), 
        .Z(n769) );
  CAOR2X1 U840 ( .A(\reg_mem[18][29] ), .B(net81941), .C(net81971), .D(n2264), 
        .Z(n770) );
  CAOR2X1 U841 ( .A(\reg_mem[18][28] ), .B(net81941), .C(net81971), .D(n2262), 
        .Z(n771) );
  CAOR2X1 U842 ( .A(\reg_mem[18][27] ), .B(net81941), .C(n1506), .D(n2260), 
        .Z(n772) );
  CAOR2X1 U843 ( .A(\reg_mem[18][26] ), .B(net81941), .C(n1506), .D(n2258), 
        .Z(n773) );
  CAOR2X1 U844 ( .A(\reg_mem[18][25] ), .B(net81941), .C(net81959), .D(n2256), 
        .Z(n774) );
  CAOR2X1 U845 ( .A(\reg_mem[18][24] ), .B(net81941), .C(net81957), .D(n2254), 
        .Z(n775) );
  CAOR2X1 U846 ( .A(\reg_mem[18][23] ), .B(n1507), .C(net81959), .D(n2252), 
        .Z(n776) );
  CAOR2X1 U847 ( .A(\reg_mem[18][22] ), .B(n1507), .C(net81957), .D(n2250), 
        .Z(n777) );
  CAOR2X1 U848 ( .A(\reg_mem[18][21] ), .B(n1507), .C(net81951), .D(n2248), 
        .Z(n778) );
  CAOR2X1 U849 ( .A(\reg_mem[18][20] ), .B(n1507), .C(net81947), .D(n2246), 
        .Z(n779) );
  CAOR2X1 U850 ( .A(\reg_mem[18][19] ), .B(n1507), .C(net81959), .D(n2244), 
        .Z(n780) );
  CAOR2X1 U851 ( .A(\reg_mem[18][18] ), .B(n1507), .C(net81957), .D(n2242), 
        .Z(n781) );
  CAOR2X1 U852 ( .A(\reg_mem[18][17] ), .B(n1507), .C(net81959), .D(n2240), 
        .Z(n782) );
  CAOR2X1 U853 ( .A(\reg_mem[18][16] ), .B(n1507), .C(net81959), .D(n2238), 
        .Z(n783) );
  CAOR2X1 U854 ( .A(\reg_mem[18][15] ), .B(n1507), .C(net81957), .D(n2236), 
        .Z(n784) );
  CAOR2X1 U855 ( .A(\reg_mem[18][14] ), .B(n1507), .C(net81957), .D(n2234), 
        .Z(n785) );
  CAOR2X1 U856 ( .A(\reg_mem[18][13] ), .B(n1507), .C(net81951), .D(net83054), 
        .Z(n786) );
  CAOR2X1 U857 ( .A(\reg_mem[18][12] ), .B(n1507), .C(net81951), .D(n2232), 
        .Z(n787) );
  CAOR2X1 U858 ( .A(\reg_mem[18][11] ), .B(n1507), .C(net81947), .D(net83058), 
        .Z(n788) );
  CAOR2X1 U859 ( .A(\reg_mem[18][10] ), .B(n1507), .C(net81945), .D(n2230), 
        .Z(n789) );
  CAOR2X1 U860 ( .A(\reg_mem[18][9] ), .B(n1507), .C(net81951), .D(n2228), .Z(
        n790) );
  CAOR2X1 U861 ( .A(\reg_mem[18][8] ), .B(n1507), .C(net81951), .D(n2226), .Z(
        n791) );
  CAOR2X1 U862 ( .A(\reg_mem[18][7] ), .B(n1507), .C(net81947), .D(n2224), .Z(
        n792) );
  CAOR2X1 U863 ( .A(\reg_mem[18][6] ), .B(n1507), .C(net81945), .D(n2222), .Z(
        n793) );
  CAOR2X1 U864 ( .A(\reg_mem[18][5] ), .B(n1507), .C(net81947), .D(n2220), .Z(
        n794) );
  CAOR2X1 U866 ( .A(\reg_mem[18][3] ), .B(n1507), .C(net81945), .D(n2218), .Z(
        n796) );
  CAOR2X1 U868 ( .A(\reg_mem[18][1] ), .B(n1507), .C(net81971), .D(n2216), .Z(
        n798) );
  CAOR2X1 U869 ( .A(\reg_mem[18][0] ), .B(n1507), .C(n1506), .D(n2214), .Z(
        n799) );
  CAOR2X1 U870 ( .A(\reg_mem[17][31] ), .B(net81981), .C(net82011), .D(n159), 
        .Z(n800) );
  CAOR2X1 U871 ( .A(\reg_mem[17][30] ), .B(net81981), .C(n1504), .D(n160), .Z(
        n801) );
  CAOR2X1 U872 ( .A(\reg_mem[17][29] ), .B(net81981), .C(net82011), .D(n161), 
        .Z(n802) );
  CAOR2X1 U873 ( .A(\reg_mem[17][28] ), .B(net81981), .C(net82011), .D(n162), 
        .Z(n803) );
  CAOR2X1 U874 ( .A(\reg_mem[17][27] ), .B(net81981), .C(n1504), .D(n163), .Z(
        n804) );
  CAOR2X1 U875 ( .A(\reg_mem[17][26] ), .B(net81981), .C(n1504), .D(n164), .Z(
        n805) );
  CAOR2X1 U876 ( .A(\reg_mem[17][25] ), .B(net81981), .C(net81999), .D(n165), 
        .Z(n806) );
  CAOR2X1 U877 ( .A(\reg_mem[17][24] ), .B(net81981), .C(net81997), .D(n166), 
        .Z(n807) );
  CAOR2X1 U878 ( .A(\reg_mem[17][23] ), .B(n1505), .C(net81999), .D(n167), .Z(
        n808) );
  CAOR2X1 U879 ( .A(\reg_mem[17][22] ), .B(n1505), .C(net81997), .D(n168), .Z(
        n809) );
  CAOR2X1 U880 ( .A(\reg_mem[17][21] ), .B(n1505), .C(net81991), .D(n169), .Z(
        n810) );
  CAOR2X1 U881 ( .A(\reg_mem[17][20] ), .B(n1505), .C(net81987), .D(n170), .Z(
        n811) );
  CAOR2X1 U882 ( .A(\reg_mem[17][19] ), .B(n1505), .C(net81999), .D(n171), .Z(
        n812) );
  CAOR2X1 U883 ( .A(\reg_mem[17][18] ), .B(n1505), .C(net81997), .D(n172), .Z(
        n813) );
  CAOR2X1 U884 ( .A(\reg_mem[17][17] ), .B(n1505), .C(net81999), .D(n173), .Z(
        n814) );
  CAOR2X1 U885 ( .A(\reg_mem[17][16] ), .B(n1505), .C(net81999), .D(n174), .Z(
        n815) );
  CAOR2X1 U886 ( .A(\reg_mem[17][15] ), .B(n1505), .C(net81997), .D(n175), .Z(
        n816) );
  CAOR2X1 U887 ( .A(\reg_mem[17][14] ), .B(n1505), .C(net81997), .D(n176), .Z(
        n817) );
  CAOR2X1 U888 ( .A(\reg_mem[17][13] ), .B(n1505), .C(net81991), .D(n177), .Z(
        n818) );
  CAOR2X1 U889 ( .A(\reg_mem[17][12] ), .B(n1505), .C(net81991), .D(n178), .Z(
        n819) );
  CAOR2X1 U890 ( .A(\reg_mem[17][11] ), .B(n1505), .C(net81987), .D(n179), .Z(
        n820) );
  CAOR2X1 U891 ( .A(\reg_mem[17][10] ), .B(n1505), .C(net81985), .D(n180), .Z(
        n821) );
  CAOR2X1 U892 ( .A(\reg_mem[17][9] ), .B(n1505), .C(net81991), .D(n181), .Z(
        n822) );
  CAOR2X1 U893 ( .A(\reg_mem[17][8] ), .B(n1505), .C(net81991), .D(n182), .Z(
        n823) );
  CAOR2X1 U894 ( .A(\reg_mem[17][7] ), .B(n1505), .C(net81987), .D(n183), .Z(
        n824) );
  CAOR2X1 U895 ( .A(\reg_mem[17][6] ), .B(n1505), .C(net81985), .D(n184), .Z(
        n825) );
  CAOR2X1 U896 ( .A(\reg_mem[17][5] ), .B(n1505), .C(net81987), .D(n185), .Z(
        n826) );
  CAOR2X1 U898 ( .A(\reg_mem[17][3] ), .B(n1505), .C(net81985), .D(n187), .Z(
        n828) );
  CAOR2X1 U900 ( .A(\reg_mem[17][1] ), .B(n1505), .C(net82011), .D(n189), .Z(
        n830) );
  CAOR2X1 U901 ( .A(\reg_mem[17][0] ), .B(n1505), .C(n1504), .D(n190), .Z(n831) );
  CAOR2X1 U902 ( .A(\reg_mem[16][31] ), .B(net82021), .C(net82051), .D(n2269), 
        .Z(n832) );
  CAOR2X1 U903 ( .A(\reg_mem[16][30] ), .B(net82021), .C(n1508), .D(n2267), 
        .Z(n833) );
  CAOR2X1 U904 ( .A(\reg_mem[16][29] ), .B(net82021), .C(net82051), .D(n2265), 
        .Z(n834) );
  CAOR2X1 U905 ( .A(\reg_mem[16][28] ), .B(net82021), .C(net82051), .D(n2263), 
        .Z(n835) );
  CAOR2X1 U906 ( .A(\reg_mem[16][27] ), .B(net82021), .C(n1508), .D(n2261), 
        .Z(n836) );
  CAOR2X1 U907 ( .A(\reg_mem[16][26] ), .B(net82021), .C(n1508), .D(n2259), 
        .Z(n837) );
  CAOR2X1 U908 ( .A(\reg_mem[16][25] ), .B(net82021), .C(net82043), .D(n2257), 
        .Z(n838) );
  CAOR2X1 U909 ( .A(\reg_mem[16][24] ), .B(net82021), .C(net82043), .D(n2255), 
        .Z(n839) );
  CAOR2X1 U910 ( .A(\reg_mem[16][23] ), .B(n1509), .C(net82039), .D(n2253), 
        .Z(n840) );
  CAOR2X1 U911 ( .A(\reg_mem[16][22] ), .B(n1509), .C(net82037), .D(n2251), 
        .Z(n841) );
  CAOR2X1 U912 ( .A(\reg_mem[16][21] ), .B(n1509), .C(net82043), .D(n2249), 
        .Z(n842) );
  CAOR2X1 U913 ( .A(\reg_mem[16][20] ), .B(n1509), .C(net82043), .D(n2247), 
        .Z(n843) );
  CAOR2X1 U914 ( .A(\reg_mem[16][19] ), .B(n1509), .C(net82039), .D(n2245), 
        .Z(n844) );
  CAOR2X1 U915 ( .A(\reg_mem[16][18] ), .B(n1509), .C(net82037), .D(n2243), 
        .Z(n845) );
  CAOR2X1 U916 ( .A(\reg_mem[16][17] ), .B(n1509), .C(net82039), .D(n2241), 
        .Z(n846) );
  CAOR2X1 U917 ( .A(\reg_mem[16][16] ), .B(n1509), .C(net82039), .D(n2239), 
        .Z(n847) );
  CAOR2X1 U918 ( .A(\reg_mem[16][15] ), .B(n1509), .C(net82037), .D(n2237), 
        .Z(n848) );
  CAOR2X1 U919 ( .A(\reg_mem[16][14] ), .B(n1509), .C(net82037), .D(n2235), 
        .Z(n849) );
  CAOR2X1 U920 ( .A(\reg_mem[16][13] ), .B(n1509), .C(net82031), .D(net83055), 
        .Z(n850) );
  CAOR2X1 U921 ( .A(\reg_mem[16][12] ), .B(n1509), .C(net82031), .D(n2233), 
        .Z(n851) );
  CAOR2X1 U922 ( .A(\reg_mem[16][11] ), .B(n1509), .C(net82027), .D(net83059), 
        .Z(n852) );
  CAOR2X1 U923 ( .A(\reg_mem[16][10] ), .B(n1509), .C(net82025), .D(n2231), 
        .Z(n853) );
  CAOR2X1 U924 ( .A(\reg_mem[16][9] ), .B(n1509), .C(net82031), .D(n2229), .Z(
        n854) );
  CAOR2X1 U925 ( .A(\reg_mem[16][8] ), .B(n1509), .C(net82031), .D(n2227), .Z(
        n855) );
  CAOR2X1 U926 ( .A(\reg_mem[16][7] ), .B(n1509), .C(net82027), .D(n2225), .Z(
        n856) );
  CAOR2X1 U927 ( .A(\reg_mem[16][6] ), .B(n1509), .C(net82025), .D(n2223), .Z(
        n857) );
  CAOR2X1 U928 ( .A(\reg_mem[16][5] ), .B(n1509), .C(net82027), .D(n2221), .Z(
        n858) );
  CAOR2X1 U930 ( .A(\reg_mem[16][3] ), .B(n1509), .C(net82025), .D(n2219), .Z(
        n860) );
  CAOR2X1 U932 ( .A(\reg_mem[16][1] ), .B(n1509), .C(net82051), .D(n2217), .Z(
        n862) );
  CAOR2X1 U933 ( .A(\reg_mem[16][0] ), .B(n1509), .C(n1508), .D(n2215), .Z(
        n863) );
  CAOR2X1 U934 ( .A(\reg_mem[15][31] ), .B(n2342), .C(n2350), .D(n2268), .Z(
        n864) );
  CAOR2X1 U935 ( .A(\reg_mem[15][30] ), .B(n2342), .C(n2349), .D(n2266), .Z(
        n865) );
  CAOR2X1 U936 ( .A(\reg_mem[15][29] ), .B(n2342), .C(n2350), .D(n2264), .Z(
        n866) );
  CAOR2X1 U937 ( .A(\reg_mem[15][28] ), .B(n2342), .C(n2350), .D(n2262), .Z(
        n867) );
  CAOR2X1 U938 ( .A(\reg_mem[15][27] ), .B(n2342), .C(n2349), .D(n2260), .Z(
        n868) );
  CAOR2X1 U939 ( .A(\reg_mem[15][26] ), .B(n2342), .C(n2349), .D(n2258), .Z(
        n869) );
  CAOR2X1 U940 ( .A(\reg_mem[15][25] ), .B(n2342), .C(n2348), .D(n2256), .Z(
        n870) );
  CAOR2X1 U941 ( .A(\reg_mem[15][24] ), .B(n2342), .C(n2348), .D(n2254), .Z(
        n871) );
  CAOR2X1 U942 ( .A(\reg_mem[15][23] ), .B(n2341), .C(n2347), .D(n2252), .Z(
        n872) );
  CAOR2X1 U943 ( .A(\reg_mem[15][22] ), .B(n2341), .C(n2346), .D(n2250), .Z(
        n873) );
  CAOR2X1 U944 ( .A(\reg_mem[15][21] ), .B(n2341), .C(n2348), .D(n2248), .Z(
        n874) );
  CAOR2X1 U945 ( .A(\reg_mem[15][20] ), .B(n2341), .C(n2348), .D(n2246), .Z(
        n875) );
  CAOR2X1 U946 ( .A(\reg_mem[15][19] ), .B(n2341), .C(n2347), .D(n2244), .Z(
        n876) );
  CAOR2X1 U947 ( .A(\reg_mem[15][18] ), .B(n2341), .C(n2346), .D(n2242), .Z(
        n877) );
  CAOR2X1 U948 ( .A(\reg_mem[15][17] ), .B(n2341), .C(n2347), .D(n2240), .Z(
        n878) );
  CAOR2X1 U949 ( .A(\reg_mem[15][16] ), .B(n2341), .C(n2347), .D(n2238), .Z(
        n879) );
  CAOR2X1 U950 ( .A(\reg_mem[15][15] ), .B(n2341), .C(n2346), .D(n2236), .Z(
        n880) );
  CAOR2X1 U951 ( .A(\reg_mem[15][14] ), .B(n2341), .C(n2346), .D(n2234), .Z(
        n881) );
  CAOR2X1 U952 ( .A(\reg_mem[15][13] ), .B(n2341), .C(n2345), .D(net83054), 
        .Z(n882) );
  CAOR2X1 U953 ( .A(\reg_mem[15][12] ), .B(n2341), .C(n2345), .D(n2232), .Z(
        n883) );
  CAOR2X1 U954 ( .A(\reg_mem[15][11] ), .B(n2340), .C(n2344), .D(net83058), 
        .Z(n884) );
  CAOR2X1 U955 ( .A(\reg_mem[15][10] ), .B(n2340), .C(n2343), .D(n2230), .Z(
        n885) );
  CAOR2X1 U956 ( .A(\reg_mem[15][9] ), .B(n2340), .C(n2345), .D(n2228), .Z(
        n886) );
  CAOR2X1 U957 ( .A(\reg_mem[15][8] ), .B(n2340), .C(n2345), .D(n2226), .Z(
        n887) );
  CAOR2X1 U958 ( .A(\reg_mem[15][7] ), .B(n2340), .C(n2344), .D(n2224), .Z(
        n888) );
  CAOR2X1 U959 ( .A(\reg_mem[15][6] ), .B(n2340), .C(n2343), .D(n2222), .Z(
        n889) );
  CAOR2X1 U960 ( .A(\reg_mem[15][5] ), .B(n2340), .C(n2344), .D(n2220), .Z(
        n890) );
  CAOR2X1 U961 ( .A(\reg_mem[15][4] ), .B(n2340), .C(n2344), .D(net83072), .Z(
        n891) );
  CAOR2X1 U962 ( .A(\reg_mem[15][3] ), .B(n2340), .C(n2343), .D(n2218), .Z(
        n892) );
  CAOR2X1 U963 ( .A(\reg_mem[15][2] ), .B(n2340), .C(n2343), .D(net83076), .Z(
        n893) );
  CAOR2X1 U964 ( .A(\reg_mem[15][1] ), .B(n2340), .C(n2350), .D(n2216), .Z(
        n894) );
  CAOR2X1 U965 ( .A(\reg_mem[15][0] ), .B(n2340), .C(n2349), .D(n2214), .Z(
        n895) );
  CAOR2X1 U966 ( .A(\reg_mem[14][31] ), .B(n2331), .C(n2338), .D(n159), .Z(
        n896) );
  CAOR2X1 U967 ( .A(\reg_mem[14][30] ), .B(n2331), .C(n2334), .D(n160), .Z(
        n897) );
  CAOR2X1 U968 ( .A(\reg_mem[14][29] ), .B(n2331), .C(n2337), .D(n161), .Z(
        n898) );
  CAOR2X1 U969 ( .A(\reg_mem[14][28] ), .B(n2331), .C(n2336), .D(n162), .Z(
        n899) );
  CAOR2X1 U970 ( .A(\reg_mem[14][27] ), .B(n2331), .C(n2333), .D(n163), .Z(
        n900) );
  CAOR2X1 U971 ( .A(\reg_mem[14][26] ), .B(n2331), .C(n2332), .D(n164), .Z(
        n901) );
  CAOR2X1 U972 ( .A(\reg_mem[14][25] ), .B(n2331), .C(n2339), .D(n165), .Z(
        n902) );
  CAOR2X1 U973 ( .A(\reg_mem[14][24] ), .B(n2331), .C(n2338), .D(n166), .Z(
        n903) );
  CAOR2X1 U974 ( .A(\reg_mem[14][23] ), .B(n1527), .C(n2339), .D(n167), .Z(
        n904) );
  CAOR2X1 U975 ( .A(\reg_mem[14][22] ), .B(n1527), .C(n2339), .D(n168), .Z(
        n905) );
  CAOR2X1 U976 ( .A(\reg_mem[14][21] ), .B(n1527), .C(n2338), .D(n169), .Z(
        n906) );
  CAOR2X1 U977 ( .A(\reg_mem[14][20] ), .B(n1527), .C(n2338), .D(n170), .Z(
        n907) );
  CAOR2X1 U978 ( .A(\reg_mem[14][19] ), .B(n1527), .C(n2337), .D(n171), .Z(
        n908) );
  CAOR2X1 U979 ( .A(\reg_mem[14][18] ), .B(n1527), .C(n2336), .D(n172), .Z(
        n909) );
  CAOR2X1 U980 ( .A(\reg_mem[14][17] ), .B(n1527), .C(n2337), .D(n173), .Z(
        n910) );
  CAOR2X1 U981 ( .A(\reg_mem[14][16] ), .B(n1527), .C(n2337), .D(n174), .Z(
        n911) );
  CAOR2X1 U982 ( .A(\reg_mem[14][15] ), .B(n1527), .C(n2336), .D(n175), .Z(
        n912) );
  CAOR2X1 U983 ( .A(\reg_mem[14][14] ), .B(n1527), .C(n2336), .D(n176), .Z(
        n913) );
  CAOR2X1 U984 ( .A(\reg_mem[14][13] ), .B(n1527), .C(n2335), .D(n177), .Z(
        n914) );
  CAOR2X1 U985 ( .A(\reg_mem[14][12] ), .B(n1527), .C(n2334), .D(n178), .Z(
        n915) );
  CAOR2X1 U986 ( .A(\reg_mem[14][11] ), .B(n1527), .C(n2335), .D(n179), .Z(
        n916) );
  CAOR2X1 U987 ( .A(\reg_mem[14][10] ), .B(n1527), .C(n2335), .D(n180), .Z(
        n917) );
  CAOR2X1 U988 ( .A(\reg_mem[14][9] ), .B(n1527), .C(n2334), .D(n181), .Z(n918) );
  CAOR2X1 U989 ( .A(\reg_mem[14][8] ), .B(n1527), .C(n2334), .D(n182), .Z(n919) );
  CAOR2X1 U990 ( .A(\reg_mem[14][7] ), .B(n1527), .C(n2333), .D(n183), .Z(n920) );
  CAOR2X1 U991 ( .A(\reg_mem[14][6] ), .B(n1527), .C(n2332), .D(n184), .Z(n921) );
  CAOR2X1 U992 ( .A(\reg_mem[14][5] ), .B(n1527), .C(n2333), .D(n185), .Z(n922) );
  CAOR2X1 U993 ( .A(\reg_mem[14][4] ), .B(n1527), .C(n2333), .D(n186), .Z(n923) );
  CAOR2X1 U994 ( .A(\reg_mem[14][3] ), .B(n220), .C(n2332), .D(n187), .Z(n924)
         );
  CAOR2X1 U995 ( .A(\reg_mem[14][2] ), .B(n220), .C(n2332), .D(n188), .Z(n925)
         );
  CAOR2X1 U996 ( .A(\reg_mem[14][1] ), .B(n220), .C(n2339), .D(n189), .Z(n926)
         );
  CAOR2X1 U997 ( .A(\reg_mem[14][0] ), .B(n220), .C(n2335), .D(n190), .Z(n927)
         );
  CAOR2X1 U998 ( .A(\reg_mem[13][31] ), .B(n2322), .C(n2330), .D(n2269), .Z(
        n928) );
  CAOR2X1 U999 ( .A(\reg_mem[13][30] ), .B(n2322), .C(n2329), .D(n2267), .Z(
        n929) );
  CAOR2X1 U1000 ( .A(\reg_mem[13][29] ), .B(n2322), .C(n2330), .D(n2265), .Z(
        n930) );
  CAOR2X1 U1001 ( .A(\reg_mem[13][28] ), .B(n2322), .C(n2330), .D(n2263), .Z(
        n931) );
  CAOR2X1 U1002 ( .A(\reg_mem[13][27] ), .B(n2322), .C(n2329), .D(n2261), .Z(
        n932) );
  CAOR2X1 U1003 ( .A(\reg_mem[13][26] ), .B(n2322), .C(n2329), .D(n2259), .Z(
        n933) );
  CAOR2X1 U1004 ( .A(\reg_mem[13][25] ), .B(n2322), .C(n2328), .D(n2257), .Z(
        n934) );
  CAOR2X1 U1005 ( .A(\reg_mem[13][24] ), .B(n2322), .C(n2328), .D(n2255), .Z(
        n935) );
  CAOR2X1 U1006 ( .A(\reg_mem[13][23] ), .B(n2321), .C(n2327), .D(n2253), .Z(
        n936) );
  CAOR2X1 U1007 ( .A(\reg_mem[13][22] ), .B(n2321), .C(n2326), .D(n2251), .Z(
        n937) );
  CAOR2X1 U1008 ( .A(\reg_mem[13][21] ), .B(n2321), .C(n2328), .D(n2249), .Z(
        n938) );
  CAOR2X1 U1009 ( .A(\reg_mem[13][20] ), .B(n2321), .C(n2328), .D(n2247), .Z(
        n939) );
  CAOR2X1 U1010 ( .A(\reg_mem[13][19] ), .B(n2321), .C(n2327), .D(n2245), .Z(
        n940) );
  CAOR2X1 U1011 ( .A(\reg_mem[13][18] ), .B(n2321), .C(n2326), .D(n2243), .Z(
        n941) );
  CAOR2X1 U1012 ( .A(\reg_mem[13][17] ), .B(n2321), .C(n2327), .D(n2241), .Z(
        n942) );
  CAOR2X1 U1013 ( .A(\reg_mem[13][16] ), .B(n2321), .C(n2327), .D(n2239), .Z(
        n943) );
  CAOR2X1 U1014 ( .A(\reg_mem[13][15] ), .B(n2321), .C(n2326), .D(n2237), .Z(
        n944) );
  CAOR2X1 U1015 ( .A(\reg_mem[13][14] ), .B(n2321), .C(n2326), .D(n2235), .Z(
        n945) );
  CAOR2X1 U1016 ( .A(\reg_mem[13][13] ), .B(n2321), .C(n2325), .D(net83055), 
        .Z(n946) );
  CAOR2X1 U1017 ( .A(\reg_mem[13][12] ), .B(n2321), .C(n2325), .D(n2233), .Z(
        n947) );
  CAOR2X1 U1018 ( .A(\reg_mem[13][11] ), .B(n2320), .C(n2324), .D(net83059), 
        .Z(n948) );
  CAOR2X1 U1019 ( .A(\reg_mem[13][10] ), .B(n2320), .C(n2323), .D(n2231), .Z(
        n949) );
  CAOR2X1 U1020 ( .A(\reg_mem[13][9] ), .B(n2320), .C(n2325), .D(n2229), .Z(
        n950) );
  CAOR2X1 U1021 ( .A(\reg_mem[13][8] ), .B(n2320), .C(n2325), .D(n2227), .Z(
        n951) );
  CAOR2X1 U1022 ( .A(\reg_mem[13][7] ), .B(n2320), .C(n2324), .D(n2225), .Z(
        n952) );
  CAOR2X1 U1023 ( .A(\reg_mem[13][6] ), .B(n2320), .C(n2323), .D(n2223), .Z(
        n953) );
  CAOR2X1 U1024 ( .A(\reg_mem[13][5] ), .B(n2320), .C(n2324), .D(n2221), .Z(
        n954) );
  CAOR2X1 U1025 ( .A(\reg_mem[13][4] ), .B(n2320), .C(n2324), .D(net83073), 
        .Z(n955) );
  CAOR2X1 U1026 ( .A(\reg_mem[13][3] ), .B(n2320), .C(n2323), .D(n2219), .Z(
        n956) );
  CAOR2X1 U1027 ( .A(\reg_mem[13][2] ), .B(n2320), .C(n2323), .D(net83077), 
        .Z(n957) );
  CAOR2X1 U1028 ( .A(\reg_mem[13][1] ), .B(n2320), .C(n2330), .D(n2217), .Z(
        n958) );
  CAOR2X1 U1029 ( .A(\reg_mem[13][0] ), .B(n2320), .C(n2329), .D(n2215), .Z(
        n959) );
  CAOR2X1 U1030 ( .A(\reg_mem[12][31] ), .B(n2311), .C(n2319), .D(n2268), .Z(
        n960) );
  CAOR2X1 U1031 ( .A(\reg_mem[12][30] ), .B(n2311), .C(n2318), .D(n2266), .Z(
        n961) );
  CAOR2X1 U1032 ( .A(\reg_mem[12][29] ), .B(n2311), .C(n2319), .D(n2264), .Z(
        n962) );
  CAOR2X1 U1033 ( .A(\reg_mem[12][28] ), .B(n2311), .C(n2319), .D(n2262), .Z(
        n963) );
  CAOR2X1 U1034 ( .A(\reg_mem[12][27] ), .B(n2311), .C(n2318), .D(n2260), .Z(
        n964) );
  CAOR2X1 U1035 ( .A(\reg_mem[12][26] ), .B(n2311), .C(n2318), .D(n2258), .Z(
        n965) );
  CAOR2X1 U1036 ( .A(\reg_mem[12][25] ), .B(n2311), .C(n2317), .D(n2256), .Z(
        n966) );
  CAOR2X1 U1037 ( .A(\reg_mem[12][24] ), .B(n2311), .C(n2317), .D(n2254), .Z(
        n967) );
  CAOR2X1 U1038 ( .A(\reg_mem[12][23] ), .B(n2310), .C(n2316), .D(n2252), .Z(
        n968) );
  CAOR2X1 U1039 ( .A(\reg_mem[12][22] ), .B(n2310), .C(n2315), .D(n2250), .Z(
        n969) );
  CAOR2X1 U1040 ( .A(\reg_mem[12][21] ), .B(n2310), .C(n2317), .D(n2248), .Z(
        n970) );
  CAOR2X1 U1041 ( .A(\reg_mem[12][20] ), .B(n2310), .C(n2317), .D(n2246), .Z(
        n971) );
  CAOR2X1 U1042 ( .A(\reg_mem[12][19] ), .B(n2310), .C(n2316), .D(n2244), .Z(
        n972) );
  CAOR2X1 U1043 ( .A(\reg_mem[12][18] ), .B(n2310), .C(n2315), .D(n2242), .Z(
        n973) );
  CAOR2X1 U1044 ( .A(\reg_mem[12][17] ), .B(n2310), .C(n2316), .D(n2240), .Z(
        n974) );
  CAOR2X1 U1045 ( .A(\reg_mem[12][16] ), .B(n2310), .C(n2316), .D(n2238), .Z(
        n975) );
  CAOR2X1 U1046 ( .A(\reg_mem[12][15] ), .B(n2310), .C(n2315), .D(n2236), .Z(
        n976) );
  CAOR2X1 U1047 ( .A(\reg_mem[12][14] ), .B(n2310), .C(n2315), .D(n2234), .Z(
        n977) );
  CAOR2X1 U1048 ( .A(\reg_mem[12][13] ), .B(n2310), .C(n2314), .D(net83054), 
        .Z(n978) );
  CAOR2X1 U1049 ( .A(\reg_mem[12][12] ), .B(n2310), .C(n2314), .D(n2232), .Z(
        n979) );
  CAOR2X1 U1050 ( .A(\reg_mem[12][11] ), .B(n2309), .C(n2313), .D(net83058), 
        .Z(n980) );
  CAOR2X1 U1051 ( .A(\reg_mem[12][10] ), .B(n2309), .C(n2312), .D(n2230), .Z(
        n981) );
  CAOR2X1 U1052 ( .A(\reg_mem[12][9] ), .B(n2309), .C(n2314), .D(n2228), .Z(
        n982) );
  CAOR2X1 U1053 ( .A(\reg_mem[12][8] ), .B(n2309), .C(n2314), .D(n2226), .Z(
        n983) );
  CAOR2X1 U1054 ( .A(\reg_mem[12][7] ), .B(n2309), .C(n2313), .D(n2224), .Z(
        n984) );
  CAOR2X1 U1055 ( .A(\reg_mem[12][6] ), .B(n2309), .C(n2312), .D(n2222), .Z(
        n985) );
  CAOR2X1 U1056 ( .A(\reg_mem[12][5] ), .B(n2309), .C(n2313), .D(n2220), .Z(
        n986) );
  CAOR2X1 U1057 ( .A(\reg_mem[12][4] ), .B(n2309), .C(n2313), .D(net83072), 
        .Z(n987) );
  CAOR2X1 U1058 ( .A(\reg_mem[12][3] ), .B(n2309), .C(n2312), .D(n2218), .Z(
        n988) );
  CAOR2X1 U1059 ( .A(\reg_mem[12][2] ), .B(n2309), .C(n2312), .D(net83076), 
        .Z(n989) );
  CAOR2X1 U1060 ( .A(\reg_mem[12][1] ), .B(n2309), .C(n2319), .D(n2216), .Z(
        n990) );
  CAOR2X1 U1061 ( .A(\reg_mem[12][0] ), .B(n2309), .C(n2318), .D(n2214), .Z(
        n991) );
  CAOR2X1 U1062 ( .A(\reg_mem[11][31] ), .B(n2304), .C(n2308), .D(n159), .Z(
        n992) );
  CAOR2X1 U1063 ( .A(\reg_mem[11][30] ), .B(n2304), .C(n2306), .D(n160), .Z(
        n993) );
  CAOR2X1 U1065 ( .A(\reg_mem[11][28] ), .B(n2304), .C(n2307), .D(n162), .Z(
        n995) );
  CAOR2X1 U1066 ( .A(\reg_mem[11][27] ), .B(n2304), .C(n2308), .D(n163), .Z(
        n996) );
  CAOR2X1 U1067 ( .A(\reg_mem[11][26] ), .B(n2304), .C(n2308), .D(n164), .Z(
        n997) );
  CAOR2X1 U1068 ( .A(\reg_mem[11][25] ), .B(n2304), .C(n2306), .D(n165), .Z(
        n998) );
  CAOR2X1 U1069 ( .A(\reg_mem[11][24] ), .B(n2304), .C(n2306), .D(n166), .Z(
        n999) );
  CAOR2X1 U1070 ( .A(\reg_mem[11][23] ), .B(n2303), .C(n2307), .D(n167), .Z(
        n1000) );
  CAOR2X1 U1071 ( .A(\reg_mem[11][22] ), .B(n2303), .C(n2307), .D(n168), .Z(
        n1001) );
  CAOR2X1 U1072 ( .A(\reg_mem[11][21] ), .B(n2303), .C(n2306), .D(n169), .Z(
        n1002) );
  CAOR2X1 U1073 ( .A(\reg_mem[11][20] ), .B(n2303), .C(n2306), .D(n170), .Z(
        n1003) );
  CAOR2X1 U1074 ( .A(\reg_mem[11][19] ), .B(n2303), .C(n2307), .D(n171), .Z(
        n1004) );
  CAOR2X1 U1075 ( .A(\reg_mem[11][18] ), .B(n2303), .C(n2307), .D(n172), .Z(
        n1005) );
  CAOR2X1 U1076 ( .A(\reg_mem[11][17] ), .B(n2303), .C(n2308), .D(n173), .Z(
        n1006) );
  CAOR2X1 U1077 ( .A(\reg_mem[11][16] ), .B(n2303), .C(n2306), .D(n174), .Z(
        n1007) );
  CAOR2X1 U1078 ( .A(\reg_mem[11][15] ), .B(n2303), .C(n2306), .D(n175), .Z(
        n1008) );
  CAOR2X1 U1079 ( .A(\reg_mem[11][14] ), .B(n2303), .C(n2306), .D(n176), .Z(
        n1009) );
  CAOR2X1 U1080 ( .A(\reg_mem[11][13] ), .B(n2303), .C(n2306), .D(n177), .Z(
        n1010) );
  CAOR2X1 U1081 ( .A(\reg_mem[11][12] ), .B(n2303), .C(n2306), .D(n178), .Z(
        n1011) );
  CAOR2X1 U1082 ( .A(\reg_mem[11][11] ), .B(n2302), .C(n2306), .D(n179), .Z(
        n1012) );
  CAOR2X1 U1083 ( .A(\reg_mem[11][10] ), .B(n2302), .C(n2306), .D(n180), .Z(
        n1013) );
  CAOR2X1 U1084 ( .A(\reg_mem[11][9] ), .B(n2302), .C(n2305), .D(n181), .Z(
        n1014) );
  CAOR2X1 U1085 ( .A(\reg_mem[11][8] ), .B(n2302), .C(n2305), .D(n182), .Z(
        n1015) );
  CAOR2X1 U1086 ( .A(\reg_mem[11][7] ), .B(n2302), .C(n2306), .D(n183), .Z(
        n1016) );
  CAOR2X1 U1087 ( .A(\reg_mem[11][6] ), .B(n2302), .C(n2306), .D(n184), .Z(
        n1017) );
  CAOR2X1 U1088 ( .A(\reg_mem[11][5] ), .B(n2302), .C(n2308), .D(n185), .Z(
        n1018) );
  CAOR2X1 U1089 ( .A(\reg_mem[11][4] ), .B(n2302), .C(n2305), .D(n186), .Z(
        n1019) );
  CAOR2X1 U1090 ( .A(\reg_mem[11][3] ), .B(n2302), .C(n2305), .D(n187), .Z(
        n1020) );
  CAOR2X1 U1091 ( .A(\reg_mem[11][2] ), .B(n2302), .C(n2307), .D(n188), .Z(
        n1021) );
  CAOR2X1 U1092 ( .A(\reg_mem[11][1] ), .B(n2302), .C(n2305), .D(n189), .Z(
        n1022) );
  CAOR2X1 U1093 ( .A(\reg_mem[11][0] ), .B(n2302), .C(n2305), .D(n190), .Z(
        n1023) );
  CAOR2X1 U1094 ( .A(\reg_mem[10][31] ), .B(n1523), .C(n2301), .D(n2269), .Z(
        n1024) );
  CAOR2X1 U1095 ( .A(\reg_mem[10][30] ), .B(n1523), .C(n2300), .D(n2267), .Z(
        n1025) );
  CAOR2X1 U1096 ( .A(\reg_mem[10][29] ), .B(n1523), .C(n2301), .D(n2265), .Z(
        n1026) );
  CAOR2X1 U1097 ( .A(\reg_mem[10][28] ), .B(n1523), .C(n2301), .D(n2263), .Z(
        n1027) );
  CAOR2X1 U1098 ( .A(\reg_mem[10][27] ), .B(n1523), .C(n2300), .D(n2261), .Z(
        n1028) );
  CAOR2X1 U1099 ( .A(\reg_mem[10][26] ), .B(n1523), .C(n2300), .D(n2259), .Z(
        n1029) );
  CAOR2X1 U1100 ( .A(\reg_mem[10][25] ), .B(n1523), .C(n2299), .D(n2257), .Z(
        n1030) );
  CAOR2X1 U1101 ( .A(\reg_mem[10][24] ), .B(n1523), .C(n2298), .D(n2255), .Z(
        n1031) );
  CAOR2X1 U1102 ( .A(\reg_mem[10][23] ), .B(n224), .C(n2299), .D(n2253), .Z(
        n1032) );
  CAOR2X1 U1103 ( .A(\reg_mem[10][22] ), .B(n224), .C(n2299), .D(n2251), .Z(
        n1033) );
  CAOR2X1 U1104 ( .A(\reg_mem[10][21] ), .B(n224), .C(n2298), .D(n2249), .Z(
        n1034) );
  CAOR2X1 U1105 ( .A(\reg_mem[10][20] ), .B(n1525), .C(n2298), .D(n2247), .Z(
        n1035) );
  CAOR2X1 U1106 ( .A(\reg_mem[10][19] ), .B(n1525), .C(n2297), .D(n2245), .Z(
        n1036) );
  CAOR2X1 U1107 ( .A(\reg_mem[10][18] ), .B(n1525), .C(n2296), .D(n2243), .Z(
        n1037) );
  CAOR2X1 U1108 ( .A(\reg_mem[10][17] ), .B(n1525), .C(n2297), .D(n2241), .Z(
        n1038) );
  CAOR2X1 U1109 ( .A(\reg_mem[10][16] ), .B(n1525), .C(n2297), .D(n2239), .Z(
        n1039) );
  CAOR2X1 U1110 ( .A(\reg_mem[10][15] ), .B(n1525), .C(n2296), .D(n2237), .Z(
        n1040) );
  CAOR2X1 U1111 ( .A(\reg_mem[10][14] ), .B(n1525), .C(n2296), .D(n2235), .Z(
        n1041) );
  CAOR2X1 U1112 ( .A(\reg_mem[10][13] ), .B(n1525), .C(n2295), .D(net83055), 
        .Z(n1042) );
  CAOR2X1 U1113 ( .A(\reg_mem[10][12] ), .B(n1525), .C(n2294), .D(n2233), .Z(
        n1043) );
  CAOR2X1 U1114 ( .A(\reg_mem[10][11] ), .B(n1525), .C(n2295), .D(net83059), 
        .Z(n1044) );
  CAOR2X1 U1115 ( .A(\reg_mem[10][10] ), .B(n1525), .C(n2295), .D(n2231), .Z(
        n1045) );
  CAOR2X1 U1116 ( .A(\reg_mem[10][9] ), .B(n1525), .C(n2294), .D(n2229), .Z(
        n1046) );
  CAOR2X1 U1117 ( .A(\reg_mem[10][8] ), .B(n1525), .C(n2294), .D(n2227), .Z(
        n1047) );
  CAOR2X1 U1118 ( .A(\reg_mem[10][7] ), .B(n1525), .C(n2293), .D(n2225), .Z(
        n1048) );
  CAOR2X1 U1119 ( .A(\reg_mem[10][6] ), .B(n1525), .C(n2293), .D(n2223), .Z(
        n1049) );
  CAOR2X1 U1120 ( .A(\reg_mem[10][5] ), .B(n1525), .C(n2292), .D(n2221), .Z(
        n1050) );
  CAOR2X1 U1121 ( .A(\reg_mem[10][4] ), .B(n1525), .C(n2292), .D(net83073), 
        .Z(n1051) );
  CAOR2X1 U1122 ( .A(\reg_mem[10][3] ), .B(n1525), .C(n1522), .D(n2219), .Z(
        n1052) );
  CAOR2X1 U1123 ( .A(\reg_mem[10][2] ), .B(n1525), .C(n1522), .D(net83077), 
        .Z(n1053) );
  CAOR2X1 U1124 ( .A(\reg_mem[10][1] ), .B(n1525), .C(n1524), .D(n2217), .Z(
        n1054) );
  CAOR2X1 U1125 ( .A(\reg_mem[10][0] ), .B(n1525), .C(n1524), .D(n2215), .Z(
        n1055) );
  CAOR2X1 U1126 ( .A(\reg_mem[9][31] ), .B(n2287), .C(n2291), .D(n2268), .Z(
        n1056) );
  CAOR2X1 U1127 ( .A(\reg_mem[9][30] ), .B(n2287), .C(n2290), .D(n2266), .Z(
        n1057) );
  CAOR2X1 U1128 ( .A(\reg_mem[9][29] ), .B(n2287), .C(n2290), .D(n2264), .Z(
        n1058) );
  CAOR2X1 U1129 ( .A(\reg_mem[9][28] ), .B(n2287), .C(n2290), .D(n2262), .Z(
        n1059) );
  CAOR2X1 U1130 ( .A(\reg_mem[9][27] ), .B(n2287), .C(n2291), .D(n2260), .Z(
        n1060) );
  CAOR2X1 U1131 ( .A(\reg_mem[9][26] ), .B(n2287), .C(n2290), .D(n2258), .Z(
        n1061) );
  CAOR2X1 U1132 ( .A(\reg_mem[9][25] ), .B(n2287), .C(n2291), .D(n2256), .Z(
        n1062) );
  CAOR2X1 U1133 ( .A(\reg_mem[9][24] ), .B(n2287), .C(n2291), .D(n2254), .Z(
        n1063) );
  CAOR2X1 U1134 ( .A(\reg_mem[9][23] ), .B(n2286), .C(n2290), .D(n2252), .Z(
        n1064) );
  CAOR2X1 U1135 ( .A(\reg_mem[9][22] ), .B(n2286), .C(n2290), .D(n2250), .Z(
        n1065) );
  CAOR2X1 U1136 ( .A(\reg_mem[9][21] ), .B(n2286), .C(n2291), .D(n2248), .Z(
        n1066) );
  CAOR2X1 U1137 ( .A(\reg_mem[9][20] ), .B(n2286), .C(n2291), .D(n2246), .Z(
        n1067) );
  CAOR2X1 U1138 ( .A(\reg_mem[9][19] ), .B(n2286), .C(n2290), .D(n2244), .Z(
        n1068) );
  CAOR2X1 U1139 ( .A(\reg_mem[9][18] ), .B(n2286), .C(n2290), .D(n2242), .Z(
        n1069) );
  CAOR2X1 U1140 ( .A(\reg_mem[9][17] ), .B(n2286), .C(n2290), .D(n2240), .Z(
        n1070) );
  CAOR2X1 U1141 ( .A(\reg_mem[9][16] ), .B(n2286), .C(n2290), .D(n2238), .Z(
        n1071) );
  CAOR2X1 U1142 ( .A(\reg_mem[9][15] ), .B(n2286), .C(n2290), .D(n2236), .Z(
        n1072) );
  CAOR2X1 U1143 ( .A(\reg_mem[9][14] ), .B(n2286), .C(n2290), .D(n2234), .Z(
        n1073) );
  CAOR2X1 U1145 ( .A(\reg_mem[9][12] ), .B(n2286), .C(n2288), .D(n2232), .Z(
        n1075) );
  CAOR2X1 U1146 ( .A(\reg_mem[9][11] ), .B(n2285), .C(n2289), .D(net83058), 
        .Z(n1076) );
  CAOR2X1 U1147 ( .A(\reg_mem[9][10] ), .B(n2285), .C(n2288), .D(n2230), .Z(
        n1077) );
  CAOR2X1 U1148 ( .A(\reg_mem[9][9] ), .B(n2285), .C(n2289), .D(n2228), .Z(
        n1078) );
  CAOR2X1 U1149 ( .A(\reg_mem[9][8] ), .B(n2285), .C(n2288), .D(n2226), .Z(
        n1079) );
  CAOR2X1 U1150 ( .A(\reg_mem[9][7] ), .B(n2285), .C(n2289), .D(n2224), .Z(
        n1080) );
  CAOR2X1 U1151 ( .A(\reg_mem[9][6] ), .B(n2285), .C(n2288), .D(n2222), .Z(
        n1081) );
  CAOR2X1 U1152 ( .A(\reg_mem[9][5] ), .B(n2285), .C(n2289), .D(n2220), .Z(
        n1082) );
  CAOR2X1 U1153 ( .A(\reg_mem[9][4] ), .B(n2285), .C(n2289), .D(net83072), .Z(
        n1083) );
  CAOR2X1 U1154 ( .A(\reg_mem[9][3] ), .B(n2285), .C(n2288), .D(n2218), .Z(
        n1084) );
  CAOR2X1 U1155 ( .A(\reg_mem[9][2] ), .B(n2285), .C(n2288), .D(net83076), .Z(
        n1085) );
  CAOR2X1 U1156 ( .A(\reg_mem[9][1] ), .B(n2285), .C(n2291), .D(n2216), .Z(
        n1086) );
  CAOR2X1 U1157 ( .A(\reg_mem[9][0] ), .B(n2285), .C(n2290), .D(n2214), .Z(
        n1087) );
  CAOR2X1 U1158 ( .A(\reg_mem[8][31] ), .B(n2280), .C(n2282), .D(n159), .Z(
        n1088) );
  CAOR2X1 U1159 ( .A(\reg_mem[8][30] ), .B(n2279), .C(n2283), .D(n160), .Z(
        n1089) );
  CAOR2X1 U1160 ( .A(\reg_mem[8][29] ), .B(n2280), .C(n2281), .D(n161), .Z(
        n1090) );
  CAOR2X1 U1161 ( .A(\reg_mem[8][28] ), .B(n2279), .C(n2283), .D(n162), .Z(
        n1091) );
  CAOR2X1 U1162 ( .A(\reg_mem[8][27] ), .B(n2279), .C(n2282), .D(n163), .Z(
        n1092) );
  CAOR2X1 U1163 ( .A(\reg_mem[8][26] ), .B(n2280), .C(n2281), .D(n164), .Z(
        n1093) );
  CAOR2X1 U1164 ( .A(\reg_mem[8][25] ), .B(n2280), .C(n2284), .D(n165), .Z(
        n1094) );
  CAOR2X1 U1165 ( .A(\reg_mem[8][24] ), .B(n2279), .C(n2284), .D(n166), .Z(
        n1095) );
  CAOR2X1 U1166 ( .A(\reg_mem[8][23] ), .B(n2280), .C(n2282), .D(n167), .Z(
        n1096) );
  CAOR2X1 U1167 ( .A(\reg_mem[8][22] ), .B(n2280), .C(n2283), .D(n168), .Z(
        n1097) );
  CAOR2X1 U1168 ( .A(\reg_mem[8][21] ), .B(n2280), .C(n2281), .D(n169), .Z(
        n1098) );
  CAOR2X1 U1169 ( .A(\reg_mem[8][20] ), .B(n2280), .C(n2283), .D(n170), .Z(
        n1099) );
  CAOR2X1 U1170 ( .A(\reg_mem[8][19] ), .B(n2280), .C(n2283), .D(n171), .Z(
        n1100) );
  CAOR2X1 U1171 ( .A(\reg_mem[8][18] ), .B(n2280), .C(n2282), .D(n172), .Z(
        n1101) );
  CAOR2X1 U1172 ( .A(\reg_mem[8][17] ), .B(n2280), .C(n2283), .D(n173), .Z(
        n1102) );
  CAOR2X1 U1173 ( .A(\reg_mem[8][16] ), .B(n2280), .C(n2283), .D(n174), .Z(
        n1103) );
  CAOR2X1 U1174 ( .A(\reg_mem[8][15] ), .B(n2280), .C(n2282), .D(n175), .Z(
        n1104) );
  CAOR2X1 U1175 ( .A(\reg_mem[8][14] ), .B(n2280), .C(n2282), .D(n176), .Z(
        n1105) );
  CAOR2X1 U1177 ( .A(\reg_mem[8][12] ), .B(n2280), .C(n2281), .D(n178), .Z(
        n1107) );
  CAOR2X1 U1178 ( .A(\reg_mem[8][11] ), .B(n2279), .C(n2282), .D(n179), .Z(
        n1108) );
  CAOR2X1 U1179 ( .A(\reg_mem[8][10] ), .B(n2279), .C(n2282), .D(n180), .Z(
        n1109) );
  CAOR2X1 U1180 ( .A(\reg_mem[8][9] ), .B(n2279), .C(n2281), .D(n181), .Z(
        n1110) );
  CAOR2X1 U1181 ( .A(\reg_mem[8][8] ), .B(n2279), .C(n2281), .D(n182), .Z(
        n1111) );
  CAOR2X1 U1182 ( .A(\reg_mem[8][7] ), .B(n2279), .C(n2283), .D(n183), .Z(
        n1112) );
  CAOR2X1 U1183 ( .A(\reg_mem[8][6] ), .B(n2279), .C(n2282), .D(n184), .Z(
        n1113) );
  CAOR2X1 U1184 ( .A(\reg_mem[8][5] ), .B(n2279), .C(n2283), .D(n185), .Z(
        n1114) );
  CAOR2X1 U1185 ( .A(\reg_mem[8][4] ), .B(n2279), .C(n2283), .D(n186), .Z(
        n1115) );
  CAOR2X1 U1186 ( .A(\reg_mem[8][3] ), .B(n2279), .C(n2281), .D(n187), .Z(
        n1116) );
  CAOR2X1 U1187 ( .A(\reg_mem[8][2] ), .B(n2279), .C(n2281), .D(n188), .Z(
        n1117) );
  CAOR2X1 U1188 ( .A(\reg_mem[8][1] ), .B(n2279), .C(n2281), .D(n189), .Z(
        n1118) );
  CAOR2X1 U1189 ( .A(\reg_mem[8][0] ), .B(n2279), .C(n2281), .D(n190), .Z(
        n1119) );
  CAOR2X1 U1190 ( .A(\reg_mem[7][31] ), .B(net82381), .C(net82403), .D(n2269), 
        .Z(n1120) );
  CAOR2X1 U1191 ( .A(\reg_mem[7][30] ), .B(net82381), .C(net82399), .D(n2267), 
        .Z(n1121) );
  CAOR2X1 U1192 ( .A(\reg_mem[7][29] ), .B(net82381), .C(net82399), .D(n2265), 
        .Z(n1122) );
  CAOR2X1 U1193 ( .A(\reg_mem[7][28] ), .B(net82381), .C(net82399), .D(n2263), 
        .Z(n1123) );
  CAOR2X1 U1194 ( .A(\reg_mem[7][27] ), .B(net82381), .C(net82403), .D(n2261), 
        .Z(n1124) );
  CAOR2X1 U1195 ( .A(\reg_mem[7][26] ), .B(net82381), .C(net82399), .D(n2259), 
        .Z(n1125) );
  CAOR2X1 U1196 ( .A(\reg_mem[7][25] ), .B(net82381), .C(net82403), .D(n2257), 
        .Z(n1126) );
  CAOR2X1 U1197 ( .A(\reg_mem[7][24] ), .B(net82381), .C(net82403), .D(n2255), 
        .Z(n1127) );
  CAOR2X1 U1198 ( .A(\reg_mem[7][23] ), .B(net82379), .C(net82399), .D(n2253), 
        .Z(n1128) );
  CAOR2X1 U1199 ( .A(\reg_mem[7][22] ), .B(net82379), .C(net82399), .D(n2251), 
        .Z(n1129) );
  CAOR2X1 U1200 ( .A(\reg_mem[7][21] ), .B(net82379), .C(net82403), .D(n2249), 
        .Z(n1130) );
  CAOR2X1 U1201 ( .A(\reg_mem[7][20] ), .B(net82379), .C(net82403), .D(n2247), 
        .Z(n1131) );
  CAOR2X1 U1202 ( .A(\reg_mem[7][19] ), .B(net82379), .C(net82399), .D(n2245), 
        .Z(n1132) );
  CAOR2X1 U1203 ( .A(\reg_mem[7][18] ), .B(net82379), .C(net82399), .D(n2243), 
        .Z(n1133) );
  CAOR2X1 U1204 ( .A(\reg_mem[7][17] ), .B(net82379), .C(net82399), .D(n2241), 
        .Z(n1134) );
  CAOR2X1 U1205 ( .A(\reg_mem[7][16] ), .B(net82379), .C(net82399), .D(n2239), 
        .Z(n1135) );
  CAOR2X1 U1206 ( .A(\reg_mem[7][15] ), .B(net82379), .C(net82399), .D(n2237), 
        .Z(n1136) );
  CAOR2X1 U1207 ( .A(\reg_mem[7][14] ), .B(net82379), .C(net82399), .D(n2235), 
        .Z(n1137) );
  CAOR2X1 U1208 ( .A(\reg_mem[7][13] ), .B(net82379), .C(net82387), .D(
        net83055), .Z(n1138) );
  CAOR2X1 U1209 ( .A(\reg_mem[7][12] ), .B(net82379), .C(net82385), .D(n2233), 
        .Z(n1139) );
  CAOR2X1 U1211 ( .A(\reg_mem[7][10] ), .B(net82377), .C(net82387), .D(n2231), 
        .Z(n1141) );
  CAOR2X1 U1212 ( .A(\reg_mem[7][9] ), .B(net82377), .C(net82387), .D(n2229), 
        .Z(n1142) );
  CAOR2X1 U1213 ( .A(\reg_mem[7][8] ), .B(net82377), .C(net82385), .D(n2227), 
        .Z(n1143) );
  CAOR2X1 U1214 ( .A(\reg_mem[7][7] ), .B(net82377), .C(net82387), .D(n2225), 
        .Z(n1144) );
  CAOR2X1 U1215 ( .A(\reg_mem[7][6] ), .B(net82377), .C(net82385), .D(n2223), 
        .Z(n1145) );
  CAOR2X1 U1216 ( .A(\reg_mem[7][5] ), .B(net82377), .C(net82387), .D(n2221), 
        .Z(n1146) );
  CAOR2X1 U1217 ( .A(\reg_mem[7][4] ), .B(net82377), .C(net82387), .D(net83073), .Z(n1147) );
  CAOR2X1 U1218 ( .A(\reg_mem[7][3] ), .B(net82377), .C(net82385), .D(n2219), 
        .Z(n1148) );
  CAOR2X1 U1219 ( .A(\reg_mem[7][2] ), .B(net82377), .C(net82385), .D(net83077), .Z(n1149) );
  CAOR2X1 U1220 ( .A(\reg_mem[7][1] ), .B(net82377), .C(net82403), .D(n2217), 
        .Z(n1150) );
  CAOR2X1 U1221 ( .A(\reg_mem[7][0] ), .B(net82377), .C(net82399), .D(n2215), 
        .Z(n1151) );
  CAOR2X1 U1222 ( .A(\reg_mem[6][31] ), .B(net82421), .C(net82437), .D(n2268), 
        .Z(n1152) );
  CAOR2X1 U1223 ( .A(\reg_mem[6][30] ), .B(net82421), .C(net82443), .D(n2266), 
        .Z(n1153) );
  CAOR2X1 U1224 ( .A(\reg_mem[6][29] ), .B(net82421), .C(net82439), .D(n2264), 
        .Z(n1154) );
  CAOR2X1 U1225 ( .A(\reg_mem[6][28] ), .B(net82421), .C(net82437), .D(n2262), 
        .Z(n1155) );
  CAOR2X1 U1226 ( .A(\reg_mem[6][27] ), .B(net82421), .C(net82443), .D(n2260), 
        .Z(n1156) );
  CAOR2X1 U1227 ( .A(\reg_mem[6][26] ), .B(net82421), .C(net82443), .D(n2258), 
        .Z(n1157) );
  CAOR2X1 U1228 ( .A(\reg_mem[6][25] ), .B(net82421), .C(net82439), .D(n2256), 
        .Z(n1158) );
  CAOR2X1 U1229 ( .A(\reg_mem[6][24] ), .B(net82421), .C(net82437), .D(n2254), 
        .Z(n1159) );
  CAOR2X1 U1230 ( .A(\reg_mem[6][23] ), .B(net82421), .C(net87043), .D(n2252), 
        .Z(n1160) );
  CAOR2X1 U1231 ( .A(\reg_mem[6][22] ), .B(net82421), .C(net82443), .D(n2250), 
        .Z(n1161) );
  CAOR2X1 U1232 ( .A(\reg_mem[6][21] ), .B(net87042), .C(net82443), .D(n2248), 
        .Z(n1162) );
  CAOR2X1 U1233 ( .A(\reg_mem[6][20] ), .B(net82421), .C(net82443), .D(n2246), 
        .Z(n1163) );
  CAOR2X1 U1234 ( .A(\reg_mem[6][19] ), .B(net87042), .C(net82439), .D(n2244), 
        .Z(n1164) );
  CAOR2X1 U1235 ( .A(\reg_mem[6][18] ), .B(net87042), .C(net82437), .D(n2242), 
        .Z(n1165) );
  CAOR2X1 U1236 ( .A(\reg_mem[6][17] ), .B(net87042), .C(net82439), .D(n2240), 
        .Z(n1166) );
  CAOR2X1 U1237 ( .A(\reg_mem[6][16] ), .B(net82421), .C(net82439), .D(n2238), 
        .Z(n1167) );
  CAOR2X1 U1238 ( .A(\reg_mem[6][15] ), .B(net87042), .C(net82437), .D(n2236), 
        .Z(n1168) );
  CAOR2X1 U1239 ( .A(\reg_mem[6][14] ), .B(n232), .C(net82437), .D(n2234), .Z(
        n1169) );
  CAOR2X1 U1240 ( .A(\reg_mem[6][13] ), .B(n232), .C(net82427), .D(net83054), 
        .Z(n1170) );
  CAOR2X1 U1241 ( .A(\reg_mem[6][12] ), .B(net87042), .C(net82425), .D(n2232), 
        .Z(n1171) );
  CAOR2X1 U1243 ( .A(\reg_mem[6][10] ), .B(n232), .C(net82427), .D(n2230), .Z(
        n1173) );
  CAOR2X1 U1244 ( .A(\reg_mem[6][9] ), .B(n232), .C(net82427), .D(n2228), .Z(
        n1174) );
  CAOR2X1 U1245 ( .A(\reg_mem[6][8] ), .B(n232), .C(net82425), .D(n2226), .Z(
        n1175) );
  CAOR2X1 U1246 ( .A(\reg_mem[6][7] ), .B(n232), .C(net82427), .D(n2224), .Z(
        n1176) );
  CAOR2X1 U1247 ( .A(\reg_mem[6][6] ), .B(n232), .C(net82425), .D(n2222), .Z(
        n1177) );
  CAOR2X1 U1248 ( .A(\reg_mem[6][5] ), .B(n232), .C(net82427), .D(n2220), .Z(
        n1178) );
  CAOR2X1 U1249 ( .A(\reg_mem[6][4] ), .B(n232), .C(net82427), .D(net83072), 
        .Z(n1179) );
  CAOR2X1 U1250 ( .A(\reg_mem[6][3] ), .B(n232), .C(net82425), .D(n2218), .Z(
        n1180) );
  CAOR2X1 U1251 ( .A(\reg_mem[6][2] ), .B(n232), .C(net82425), .D(net83076), 
        .Z(n1181) );
  CAOR2X1 U1252 ( .A(\reg_mem[6][1] ), .B(n232), .C(net82439), .D(n2216), .Z(
        n1182) );
  CAOR2X1 U1253 ( .A(\reg_mem[6][0] ), .B(n232), .C(net82443), .D(n2214), .Z(
        n1183) );
  CAOR2X1 U1254 ( .A(\reg_mem[5][31] ), .B(net82461), .C(net82491), .D(n159), 
        .Z(n1184) );
  CAOR2X1 U1255 ( .A(\reg_mem[5][30] ), .B(net82461), .C(net82489), .D(n160), 
        .Z(n1185) );
  CAOR2X1 U1256 ( .A(\reg_mem[5][29] ), .B(net82461), .C(net82491), .D(n161), 
        .Z(n1186) );
  CAOR2X1 U1257 ( .A(\reg_mem[5][28] ), .B(net82461), .C(net82491), .D(n162), 
        .Z(n1187) );
  CAOR2X1 U1258 ( .A(\reg_mem[5][27] ), .B(net82461), .C(net82489), .D(n163), 
        .Z(n1188) );
  CAOR2X1 U1259 ( .A(\reg_mem[5][26] ), .B(net82461), .C(net82489), .D(n164), 
        .Z(n1189) );
  CAOR2X1 U1260 ( .A(\reg_mem[5][25] ), .B(net82461), .C(net82485), .D(n165), 
        .Z(n1190) );
  CAOR2X1 U1261 ( .A(\reg_mem[5][24] ), .B(net82461), .C(net82483), .D(n166), 
        .Z(n1191) );
  CAOR2X1 U1262 ( .A(\reg_mem[5][23] ), .B(net82459), .C(net82485), .D(n167), 
        .Z(n1192) );
  CAOR2X1 U1263 ( .A(\reg_mem[5][22] ), .B(net82459), .C(net82485), .D(n168), 
        .Z(n1193) );
  CAOR2X1 U1264 ( .A(\reg_mem[5][21] ), .B(net82459), .C(net82483), .D(n169), 
        .Z(n1194) );
  CAOR2X1 U1265 ( .A(\reg_mem[5][20] ), .B(net82459), .C(net82483), .D(n170), 
        .Z(n1195) );
  CAOR2X1 U1266 ( .A(\reg_mem[5][19] ), .B(net82459), .C(net82479), .D(n171), 
        .Z(n1196) );
  CAOR2X1 U1267 ( .A(\reg_mem[5][18] ), .B(net82459), .C(net82477), .D(n172), 
        .Z(n1197) );
  CAOR2X1 U1268 ( .A(\reg_mem[5][17] ), .B(net82459), .C(net82479), .D(n173), 
        .Z(n1198) );
  CAOR2X1 U1269 ( .A(\reg_mem[5][16] ), .B(net82459), .C(net82479), .D(n174), 
        .Z(n1199) );
  CAOR2X1 U1270 ( .A(\reg_mem[5][15] ), .B(net82459), .C(net82477), .D(n175), 
        .Z(n1200) );
  CAOR2X1 U1271 ( .A(\reg_mem[5][14] ), .B(net82459), .C(net82477), .D(n176), 
        .Z(n1201) );
  CAOR2X1 U1272 ( .A(\reg_mem[5][13] ), .B(net82459), .C(net82473), .D(n177), 
        .Z(n1202) );
  CAOR2X1 U1273 ( .A(\reg_mem[5][12] ), .B(net82459), .C(net82469), .D(n178), 
        .Z(n1203) );
  CAOR2X1 U1275 ( .A(\reg_mem[5][10] ), .B(net82457), .C(net82473), .D(n180), 
        .Z(n1205) );
  CAOR2X1 U1276 ( .A(\reg_mem[5][9] ), .B(net82457), .C(net82489), .D(n181), 
        .Z(n1206) );
  CAOR2X1 U1278 ( .A(\reg_mem[5][7] ), .B(net82457), .C(net82469), .D(n183), 
        .Z(n1208) );
  CAOR2X1 U1279 ( .A(\reg_mem[5][6] ), .B(net82457), .C(net82469), .D(n184), 
        .Z(n1209) );
  CAOR2X1 U1280 ( .A(\reg_mem[5][5] ), .B(net82457), .C(net82465), .D(n185), 
        .Z(n1210) );
  CAOR2X1 U1281 ( .A(\reg_mem[5][4] ), .B(net82457), .C(net82463), .D(n186), 
        .Z(n1211) );
  CAOR2X1 U1282 ( .A(\reg_mem[5][3] ), .B(net82457), .C(net82465), .D(n187), 
        .Z(n1212) );
  CAOR2X1 U1283 ( .A(\reg_mem[5][2] ), .B(net82457), .C(net82465), .D(n188), 
        .Z(n1213) );
  CAOR2X1 U1284 ( .A(\reg_mem[5][1] ), .B(net82457), .C(net82463), .D(n189), 
        .Z(n1214) );
  CAOR2X1 U1285 ( .A(\reg_mem[5][0] ), .B(net82457), .C(net82463), .D(n190), 
        .Z(n1215) );
  CAOR2X1 U1286 ( .A(\reg_mem[4][31] ), .B(net82501), .C(net82533), .D(n2269), 
        .Z(n1216) );
  CAOR2X1 U1287 ( .A(\reg_mem[4][30] ), .B(net82501), .C(net82533), .D(n2267), 
        .Z(n1217) );
  CAOR2X1 U1288 ( .A(\reg_mem[4][29] ), .B(net82501), .C(net82529), .D(n2265), 
        .Z(n1218) );
  CAOR2X1 U1289 ( .A(\reg_mem[4][28] ), .B(net82501), .C(net82527), .D(n2263), 
        .Z(n1219) );
  CAOR2X1 U1290 ( .A(\reg_mem[4][27] ), .B(net82501), .C(net82529), .D(n2261), 
        .Z(n1220) );
  CAOR2X1 U1291 ( .A(\reg_mem[4][26] ), .B(net82501), .C(net82529), .D(n2259), 
        .Z(n1221) );
  CAOR2X1 U1292 ( .A(\reg_mem[4][25] ), .B(net82501), .C(net82527), .D(n2257), 
        .Z(n1222) );
  CAOR2X1 U1293 ( .A(\reg_mem[4][24] ), .B(net82501), .C(net82527), .D(n2255), 
        .Z(n1223) );
  CAOR2X1 U1294 ( .A(\reg_mem[4][23] ), .B(net82499), .C(net82523), .D(n2253), 
        .Z(n1224) );
  CAOR2X1 U1295 ( .A(\reg_mem[4][22] ), .B(net82499), .C(net82521), .D(n2251), 
        .Z(n1225) );
  CAOR2X1 U1296 ( .A(\reg_mem[4][21] ), .B(net82499), .C(net82523), .D(n2249), 
        .Z(n1226) );
  CAOR2X1 U1297 ( .A(\reg_mem[4][20] ), .B(net82499), .C(net82523), .D(n2247), 
        .Z(n1227) );
  CAOR2X1 U1298 ( .A(\reg_mem[4][19] ), .B(net82499), .C(net82521), .D(n2245), 
        .Z(n1228) );
  CAOR2X1 U1299 ( .A(\reg_mem[4][18] ), .B(net82499), .C(net82521), .D(n2243), 
        .Z(n1229) );
  CAOR2X1 U1300 ( .A(\reg_mem[4][17] ), .B(net82499), .C(net82519), .D(n2241), 
        .Z(n1230) );
  CAOR2X1 U1301 ( .A(\reg_mem[4][16] ), .B(net82499), .C(net82519), .D(n2239), 
        .Z(n1231) );
  CAOR2X1 U1302 ( .A(\reg_mem[4][15] ), .B(net82499), .C(net82517), .D(n2237), 
        .Z(n1232) );
  CAOR2X1 U1303 ( .A(\reg_mem[4][14] ), .B(net82499), .C(net82517), .D(n2235), 
        .Z(n1233) );
  CAOR2X1 U1304 ( .A(\reg_mem[4][13] ), .B(net82499), .C(net82515), .D(
        net83055), .Z(n1234) );
  CAOR2X1 U1305 ( .A(\reg_mem[4][12] ), .B(net82499), .C(net82515), .D(n2233), 
        .Z(n1235) );
  CAOR2X1 U1307 ( .A(\reg_mem[4][10] ), .B(net82497), .C(net82513), .D(n2231), 
        .Z(n1237) );
  CAOR2X1 U1308 ( .A(\reg_mem[4][9] ), .B(net82497), .C(net82533), .D(n2229), 
        .Z(n1238) );
  CAOR2X1 U1310 ( .A(\reg_mem[4][7] ), .B(net82497), .C(net82509), .D(n2225), 
        .Z(n1240) );
  CAOR2X1 U1311 ( .A(\reg_mem[4][6] ), .B(net82497), .C(net82509), .D(n2223), 
        .Z(n1241) );
  CAOR2X1 U1312 ( .A(\reg_mem[4][5] ), .B(net82497), .C(net82507), .D(n2221), 
        .Z(n1242) );
  CAOR2X1 U1313 ( .A(\reg_mem[4][4] ), .B(net82497), .C(net82507), .D(net83073), .Z(n1243) );
  CAOR2X1 U1314 ( .A(\reg_mem[4][3] ), .B(net82497), .C(net82505), .D(n2219), 
        .Z(n1244) );
  CAOR2X1 U1315 ( .A(\reg_mem[4][2] ), .B(net82497), .C(net82505), .D(net83077), .Z(n1245) );
  CAOR2X1 U1316 ( .A(\reg_mem[4][1] ), .B(net82497), .C(net82503), .D(n2217), 
        .Z(n1246) );
  CAOR2X1 U1317 ( .A(\reg_mem[4][0] ), .B(net82497), .C(net82503), .D(n2215), 
        .Z(n1247) );
  CAOR2X1 U1318 ( .A(\reg_mem[3][31] ), .B(net82541), .C(net82571), .D(n2268), 
        .Z(n1248) );
  CAOR2X1 U1319 ( .A(\reg_mem[3][30] ), .B(net82541), .C(net82557), .D(n2266), 
        .Z(n1249) );
  CAOR2X1 U1320 ( .A(\reg_mem[3][29] ), .B(net82541), .C(net82571), .D(n2264), 
        .Z(n1250) );
  CAOR2X1 U1321 ( .A(\reg_mem[3][28] ), .B(net82541), .C(net82571), .D(n2262), 
        .Z(n1251) );
  CAOR2X1 U1322 ( .A(\reg_mem[3][27] ), .B(net82541), .C(net82557), .D(n2260), 
        .Z(n1252) );
  CAOR2X1 U1323 ( .A(\reg_mem[3][26] ), .B(net82541), .C(net82549), .D(n2258), 
        .Z(n1253) );
  CAOR2X1 U1324 ( .A(\reg_mem[3][25] ), .B(net82541), .C(net82549), .D(n2256), 
        .Z(n1254) );
  CAOR2X1 U1325 ( .A(\reg_mem[3][24] ), .B(net82541), .C(net82549), .D(n2254), 
        .Z(n1255) );
  CAOR2X1 U1326 ( .A(\reg_mem[3][23] ), .B(net82539), .C(net82549), .D(n2252), 
        .Z(n1256) );
  CAOR2X1 U1327 ( .A(\reg_mem[3][22] ), .B(net82539), .C(net82557), .D(n2250), 
        .Z(n1257) );
  CAOR2X1 U1328 ( .A(\reg_mem[3][21] ), .B(net82539), .C(net82549), .D(n2248), 
        .Z(n1258) );
  CAOR2X1 U1329 ( .A(\reg_mem[3][20] ), .B(net82539), .C(net82549), .D(n2246), 
        .Z(n1259) );
  CAOR2X1 U1330 ( .A(\reg_mem[3][19] ), .B(net82539), .C(net82571), .D(n2244), 
        .Z(n1260) );
  CAOR2X1 U1331 ( .A(\reg_mem[3][18] ), .B(net82539), .C(net82557), .D(n2242), 
        .Z(n1261) );
  CAOR2X1 U1332 ( .A(\reg_mem[3][17] ), .B(net82539), .C(net82557), .D(n2240), 
        .Z(n1262) );
  CAOR2X1 U1333 ( .A(\reg_mem[3][16] ), .B(net82539), .C(net82549), .D(n2238), 
        .Z(n1263) );
  CAOR2X1 U1334 ( .A(\reg_mem[3][15] ), .B(net82539), .C(net82557), .D(n2236), 
        .Z(n1264) );
  CAOR2X1 U1335 ( .A(\reg_mem[3][14] ), .B(net82539), .C(net82557), .D(n2234), 
        .Z(n1265) );
  CAOR2X1 U1337 ( .A(\reg_mem[3][12] ), .B(net82539), .C(net82549), .D(n2232), 
        .Z(n1267) );
  CAOR2X1 U1338 ( .A(\reg_mem[3][11] ), .B(net82537), .C(net82543), .D(
        net83058), .Z(n1268) );
  CAOR2X1 U1339 ( .A(\reg_mem[3][10] ), .B(net82537), .C(net82543), .D(n2230), 
        .Z(n1269) );
  CAOR2X1 U1340 ( .A(\reg_mem[3][9] ), .B(net82537), .C(net82549), .D(n2228), 
        .Z(n1270) );
  CAOR2X1 U1342 ( .A(\reg_mem[3][7] ), .B(net82537), .C(net82549), .D(n2224), 
        .Z(n1272) );
  CAOR2X1 U1343 ( .A(\reg_mem[3][6] ), .B(net82537), .C(net82549), .D(n2222), 
        .Z(n1273) );
  CAOR2X1 U1344 ( .A(\reg_mem[3][5] ), .B(net82537), .C(net82571), .D(n2220), 
        .Z(n1274) );
  CAOR2X1 U1345 ( .A(\reg_mem[3][4] ), .B(net82537), .C(net82543), .D(net83072), .Z(n1275) );
  CAOR2X1 U1346 ( .A(\reg_mem[3][3] ), .B(net82537), .C(net82543), .D(n2218), 
        .Z(n1276) );
  CAOR2X1 U1347 ( .A(\reg_mem[3][2] ), .B(net82537), .C(net82549), .D(net83076), .Z(n1277) );
  CAOR2X1 U1348 ( .A(\reg_mem[3][1] ), .B(net82537), .C(net82543), .D(n2216), 
        .Z(n1278) );
  CAOR2X1 U1349 ( .A(\reg_mem[3][0] ), .B(net82537), .C(net82543), .D(n2214), 
        .Z(n1279) );
  CAOR2X1 U1350 ( .A(\reg_mem[2][31] ), .B(net82581), .C(net82611), .D(n159), 
        .Z(n1280) );
  CAOR2X1 U1351 ( .A(\reg_mem[2][30] ), .B(net82581), .C(net82609), .D(n160), 
        .Z(n1281) );
  CAOR2X1 U1352 ( .A(\reg_mem[2][29] ), .B(net82581), .C(net82611), .D(n161), 
        .Z(n1282) );
  CAOR2X1 U1353 ( .A(\reg_mem[2][28] ), .B(net82581), .C(net82611), .D(n162), 
        .Z(n1283) );
  CAOR2X1 U1354 ( .A(\reg_mem[2][27] ), .B(net82581), .C(net82609), .D(n163), 
        .Z(n1284) );
  CAOR2X1 U1355 ( .A(\reg_mem[2][26] ), .B(net82581), .C(net82609), .D(n164), 
        .Z(n1285) );
  CAOR2X1 U1356 ( .A(\reg_mem[2][25] ), .B(net82581), .C(net82605), .D(n165), 
        .Z(n1286) );
  CAOR2X1 U1357 ( .A(\reg_mem[2][24] ), .B(net82581), .C(net82603), .D(n166), 
        .Z(n1287) );
  CAOR2X1 U1358 ( .A(\reg_mem[2][23] ), .B(net82579), .C(net82605), .D(n167), 
        .Z(n1288) );
  CAOR2X1 U1359 ( .A(\reg_mem[2][22] ), .B(net82579), .C(net82605), .D(n168), 
        .Z(n1289) );
  CAOR2X1 U1360 ( .A(\reg_mem[2][21] ), .B(net82579), .C(net82603), .D(n169), 
        .Z(n1290) );
  CAOR2X1 U1361 ( .A(\reg_mem[2][20] ), .B(net82579), .C(net82603), .D(n170), 
        .Z(n1291) );
  CAOR2X1 U1362 ( .A(\reg_mem[2][19] ), .B(net82579), .C(net82599), .D(n171), 
        .Z(n1292) );
  CAOR2X1 U1363 ( .A(\reg_mem[2][18] ), .B(net82579), .C(net82597), .D(n172), 
        .Z(n1293) );
  CAOR2X1 U1364 ( .A(\reg_mem[2][17] ), .B(net82579), .C(net82599), .D(n173), 
        .Z(n1294) );
  CAOR2X1 U1365 ( .A(\reg_mem[2][16] ), .B(net82579), .C(net82599), .D(n174), 
        .Z(n1295) );
  CAOR2X1 U1366 ( .A(\reg_mem[2][15] ), .B(net82579), .C(net82597), .D(n175), 
        .Z(n1296) );
  CAOR2X1 U1367 ( .A(\reg_mem[2][14] ), .B(net82579), .C(net82597), .D(n176), 
        .Z(n1297) );
  CAOR2X1 U1369 ( .A(\reg_mem[2][12] ), .B(net82579), .C(net82593), .D(n178), 
        .Z(n1299) );
  CAOR2X1 U1370 ( .A(\reg_mem[2][11] ), .B(net82577), .C(net82593), .D(n179), 
        .Z(n1300) );
  CAOR2X1 U1371 ( .A(\reg_mem[2][10] ), .B(net82577), .C(net82593), .D(n180), 
        .Z(n1301) );
  CAOR2X1 U1372 ( .A(\reg_mem[2][9] ), .B(net82577), .C(net82591), .D(n181), 
        .Z(n1302) );
  CAOR2X1 U1373 ( .A(\reg_mem[2][8] ), .B(net82577), .C(net82591), .D(n182), 
        .Z(n1303) );
  CAOR2X1 U1374 ( .A(\reg_mem[2][7] ), .B(net82577), .C(net82587), .D(n183), 
        .Z(n1304) );
  CAOR2X1 U1375 ( .A(\reg_mem[2][6] ), .B(net82577), .C(net82585), .D(n184), 
        .Z(n1305) );
  CAOR2X1 U1376 ( .A(\reg_mem[2][5] ), .B(net82577), .C(net82587), .D(n185), 
        .Z(n1306) );
  CAOR2X1 U1377 ( .A(\reg_mem[2][4] ), .B(net82577), .C(net82587), .D(n186), 
        .Z(n1307) );
  CAOR2X1 U1378 ( .A(\reg_mem[2][3] ), .B(net82577), .C(net82585), .D(n187), 
        .Z(n1308) );
  CAOR2X1 U1379 ( .A(\reg_mem[2][2] ), .B(net82577), .C(net82585), .D(n188), 
        .Z(n1309) );
  CAOR2X1 U1380 ( .A(\reg_mem[2][1] ), .B(net82577), .C(net82583), .D(n189), 
        .Z(n1310) );
  CAOR2X1 U1381 ( .A(\reg_mem[2][0] ), .B(net82577), .C(net82583), .D(n190), 
        .Z(n1311) );
  CAOR2X1 U1382 ( .A(\reg_mem[1][31] ), .B(net82621), .C(net82643), .D(n2269), 
        .Z(n1312) );
  CAOR2X1 U1383 ( .A(\reg_mem[1][30] ), .B(net82621), .C(net82639), .D(n2267), 
        .Z(n1313) );
  CAOR2X1 U1384 ( .A(\reg_mem[1][29] ), .B(net82621), .C(net82639), .D(n2265), 
        .Z(n1314) );
  CAOR2X1 U1385 ( .A(\reg_mem[1][28] ), .B(net82621), .C(net82639), .D(n2263), 
        .Z(n1315) );
  CAOR2X1 U1386 ( .A(\reg_mem[1][27] ), .B(net82621), .C(net82643), .D(n2261), 
        .Z(n1316) );
  CAOR2X1 U1387 ( .A(\reg_mem[1][26] ), .B(net82621), .C(net82639), .D(n2259), 
        .Z(n1317) );
  CAOR2X1 U1388 ( .A(\reg_mem[1][25] ), .B(net82621), .C(net82643), .D(n2257), 
        .Z(n1318) );
  CAOR2X1 U1389 ( .A(\reg_mem[1][24] ), .B(net82621), .C(net82643), .D(n2255), 
        .Z(n1319) );
  CAOR2X1 U1390 ( .A(\reg_mem[1][23] ), .B(net82619), .C(net82639), .D(n2253), 
        .Z(n1320) );
  CAOR2X1 U1391 ( .A(\reg_mem[1][22] ), .B(net82619), .C(net82639), .D(n2251), 
        .Z(n1321) );
  CAOR2X1 U1392 ( .A(\reg_mem[1][21] ), .B(net82619), .C(net82643), .D(n2249), 
        .Z(n1322) );
  CAOR2X1 U1393 ( .A(\reg_mem[1][20] ), .B(net82619), .C(net82643), .D(n2247), 
        .Z(n1323) );
  CAOR2X1 U1394 ( .A(\reg_mem[1][19] ), .B(net82619), .C(net82639), .D(n2245), 
        .Z(n1324) );
  CAOR2X1 U1395 ( .A(\reg_mem[1][18] ), .B(net82619), .C(net82639), .D(n2243), 
        .Z(n1325) );
  CAOR2X1 U1396 ( .A(\reg_mem[1][17] ), .B(net82619), .C(net82639), .D(n2241), 
        .Z(n1326) );
  CAOR2X1 U1397 ( .A(\reg_mem[1][16] ), .B(net82619), .C(net82639), .D(n2239), 
        .Z(n1327) );
  CAOR2X1 U1398 ( .A(\reg_mem[1][15] ), .B(net82619), .C(net82639), .D(n2237), 
        .Z(n1328) );
  CAOR2X1 U1399 ( .A(\reg_mem[1][14] ), .B(net82619), .C(net82639), .D(n2235), 
        .Z(n1329) );
  CAOR2X1 U1401 ( .A(\reg_mem[1][12] ), .B(net82619), .C(net82627), .D(n2233), 
        .Z(n1331) );
  CAOR2X1 U1402 ( .A(\reg_mem[1][11] ), .B(net82617), .C(net82627), .D(
        net83059), .Z(n1332) );
  CAOR2X1 U1403 ( .A(\reg_mem[1][10] ), .B(net82617), .C(net82625), .D(n2231), 
        .Z(n1333) );
  CAOR2X1 U1404 ( .A(\reg_mem[1][9] ), .B(net82617), .C(net82627), .D(n2229), 
        .Z(n1334) );
  CAOR2X1 U1405 ( .A(\reg_mem[1][8] ), .B(net82617), .C(net82625), .D(n2227), 
        .Z(n1335) );
  CAOR2X1 U1406 ( .A(\reg_mem[1][7] ), .B(net82617), .C(net82627), .D(n2225), 
        .Z(n1336) );
  CAOR2X1 U1407 ( .A(\reg_mem[1][6] ), .B(net82617), .C(net82625), .D(n2223), 
        .Z(n1337) );
  CAOR2X1 U1408 ( .A(\reg_mem[1][5] ), .B(net82617), .C(net82627), .D(n2221), 
        .Z(n1338) );
  CAOR2X1 U1409 ( .A(\reg_mem[1][4] ), .B(net82617), .C(net82627), .D(net83073), .Z(n1339) );
  CAOR2X1 U1410 ( .A(\reg_mem[1][3] ), .B(net82617), .C(net82625), .D(n2219), 
        .Z(n1340) );
  CAOR2X1 U1411 ( .A(\reg_mem[1][2] ), .B(net82617), .C(net82625), .D(net83077), .Z(n1341) );
  CAOR2X1 U1412 ( .A(\reg_mem[1][1] ), .B(net82617), .C(net82643), .D(n2217), 
        .Z(n1342) );
  CAOR2X1 U1413 ( .A(\reg_mem[1][0] ), .B(net82617), .C(net82639), .D(n2215), 
        .Z(n1343) );
  CAOR2X1 U1414 ( .A(\reg_mem[0][31] ), .B(n1530), .C(net82683), .D(n2268), 
        .Z(n1344) );
  CAOR2X1 U1415 ( .A(data_mem_rdata_i[31]), .B(n2202), .C(alu_op_wb[31]), .D(
        n2211), .Z(n159) );
  CAOR2X1 U1416 ( .A(\reg_mem[0][30] ), .B(n1530), .C(net82689), .D(n2266), 
        .Z(n1345) );
  CAOR2X1 U1418 ( .A(\reg_mem[0][29] ), .B(n1530), .C(net82679), .D(n2264), 
        .Z(n1346) );
  CAOR2X1 U1420 ( .A(\reg_mem[0][28] ), .B(n1530), .C(net82677), .D(n2262), 
        .Z(n1347) );
  CAOR2X1 U1422 ( .A(\reg_mem[0][27] ), .B(n1530), .C(net82689), .D(n2260), 
        .Z(n1348) );
  CAOR2X1 U1424 ( .A(\reg_mem[0][26] ), .B(n1530), .C(net82689), .D(n2258), 
        .Z(n1349) );
  CAOR2X1 U1426 ( .A(\reg_mem[0][25] ), .B(n1530), .C(net82683), .D(n2256), 
        .Z(n1350) );
  CAOR2X1 U1428 ( .A(\reg_mem[0][24] ), .B(n1530), .C(net82683), .D(n2254), 
        .Z(n1351) );
  CAOR2X1 U1430 ( .A(\reg_mem[0][23] ), .B(n1530), .C(net82679), .D(n2252), 
        .Z(n1352) );
  CAOR2X1 U1432 ( .A(\reg_mem[0][22] ), .B(n1530), .C(net82677), .D(n2250), 
        .Z(n1353) );
  CAOR2X1 U1434 ( .A(\reg_mem[0][21] ), .B(n1530), .C(net82683), .D(n2248), 
        .Z(n1354) );
  CAOR2X1 U1436 ( .A(\reg_mem[0][20] ), .B(n1530), .C(net82683), .D(n2246), 
        .Z(n1355) );
  CAOR2X1 U1438 ( .A(\reg_mem[0][19] ), .B(n1530), .C(net82679), .D(n2244), 
        .Z(n1356) );
  CAOR2X1 U1440 ( .A(\reg_mem[0][18] ), .B(n1530), .C(net82677), .D(n2242), 
        .Z(n1357) );
  CAOR2X1 U1442 ( .A(\reg_mem[0][17] ), .B(n1530), .C(net82679), .D(n2240), 
        .Z(n1358) );
  CAOR2X1 U1444 ( .A(\reg_mem[0][16] ), .B(n1530), .C(net82679), .D(n2238), 
        .Z(n1359) );
  CAOR2X1 U1446 ( .A(\reg_mem[0][15] ), .B(n1530), .C(net82677), .D(n2236), 
        .Z(n1360) );
  CAOR2X1 U1448 ( .A(\reg_mem[0][14] ), .B(n238), .C(net82677), .D(n2234), .Z(
        n1361) );
  CAOR2X1 U1452 ( .A(\reg_mem[0][12] ), .B(n238), .C(net82667), .D(n2232), .Z(
        n1363) );
  CAOR2X1 U1453 ( .A(data_mem_rdata_i[12]), .B(n2202), .C(alu_op_wb[12]), .D(
        n2210), .Z(n178) );
  CAOR2X1 U1454 ( .A(\reg_mem[0][11] ), .B(n238), .C(net82667), .D(net83058), 
        .Z(n1364) );
  CAOR2X1 U1455 ( .A(data_mem_rdata_i[11]), .B(n2202), .C(alu_op_wb[11]), .D(
        n2209), .Z(n179) );
  CAOR2X1 U1456 ( .A(\reg_mem[0][10] ), .B(n238), .C(net82665), .D(n2230), .Z(
        n1365) );
  CAOR2X1 U1457 ( .A(data_mem_rdata_i[10]), .B(n2202), .C(alu_op_wb[10]), .D(
        n2208), .Z(n180) );
  CAOR2X1 U1458 ( .A(\reg_mem[0][9] ), .B(n238), .C(net82667), .D(n2228), .Z(
        n1366) );
  CAOR2X1 U1459 ( .A(data_mem_rdata_i[9]), .B(n2202), .C(alu_op_wb[9]), .D(
        n2206), .Z(n181) );
  CAOR2X1 U1460 ( .A(\reg_mem[0][8] ), .B(n238), .C(net82665), .D(n2226), .Z(
        n1367) );
  CAOR2X1 U1461 ( .A(data_mem_rdata_i[8]), .B(n2202), .C(alu_op_wb[8]), .D(
        n2205), .Z(n182) );
  CAOR2X1 U1462 ( .A(\reg_mem[0][7] ), .B(n238), .C(net82667), .D(n2224), .Z(
        n1368) );
  CAOR2X1 U1463 ( .A(data_mem_rdata_i[7]), .B(n2202), .C(alu_op_wb[7]), .D(
        n2204), .Z(n183) );
  CAOR2X1 U1464 ( .A(\reg_mem[0][6] ), .B(n238), .C(net82665), .D(n2222), .Z(
        n1369) );
  CAOR2X1 U1465 ( .A(data_mem_rdata_i[6]), .B(n2202), .C(alu_op_wb[6]), .D(
        n2204), .Z(n184) );
  CAOR2X1 U1466 ( .A(\reg_mem[0][5] ), .B(n238), .C(net82667), .D(n2220), .Z(
        n1370) );
  CAOR2X1 U1467 ( .A(data_mem_rdata_i[5]), .B(n2202), .C(alu_op_wb[5]), .D(
        n2205), .Z(n185) );
  CAOR2X1 U1468 ( .A(\reg_mem[0][4] ), .B(n238), .C(net82667), .D(net83072), 
        .Z(n1371) );
  CAOR2X1 U1469 ( .A(data_mem_rdata_i[4]), .B(n2202), .C(alu_op_wb[4]), .D(
        n2204), .Z(n186) );
  CAOR2X1 U1470 ( .A(\reg_mem[0][3] ), .B(n1530), .C(net82665), .D(n2218), .Z(
        n1372) );
  CAOR2X1 U1471 ( .A(data_mem_rdata_i[3]), .B(n2202), .C(alu_op_wb[3]), .D(
        n2207), .Z(n187) );
  CAOR2X1 U1472 ( .A(\reg_mem[0][2] ), .B(n1530), .C(net82665), .D(net83076), 
        .Z(n1373) );
  CAOR2X1 U1473 ( .A(data_mem_rdata_i[2]), .B(n2202), .C(alu_op_wb[2]), .D(
        n2206), .Z(n188) );
  CAOR2X1 U1474 ( .A(\reg_mem[0][1] ), .B(n1530), .C(net82689), .D(n2216), .Z(
        n1374) );
  CAOR2X1 U1475 ( .A(data_mem_rdata_i[1]), .B(n2202), .C(alu_op_wb[1]), .D(
        n2205), .Z(n189) );
  CAOR2X1 U1476 ( .A(\reg_mem[0][0] ), .B(n1530), .C(net82689), .D(n2214), .Z(
        n1375) );
  CAOR2X1 U1477 ( .A(data_mem_rdata_i[0]), .B(n2202), .C(alu_op_wb[0]), .D(
        n2204), .Z(n190) );
  COR2X1 U1478 ( .A(data_mem_rd_d), .B(i_type_wb), .Z(n241) );
  COR2X1 U1479 ( .A(i_type_wb), .B(n240), .Z(n239) );
  COR2X1 U1480 ( .A(j_type_wb), .B(r_type_wb), .Z(n240) );
  CAN4X1 U1488 ( .A(n99), .B(n98), .C(n100), .D(n248), .Z(n243) );
  CFD2QX2 \regA_reg[31]  ( .D(N300), .CP(clk), .CD(rst), .Q(regA[31]) );
  CFD2QX2 \regA_reg[30]  ( .D(N299), .CP(clk), .CD(rst), .Q(regA[30]) );
  CFD2QX2 \regA_reg[2]  ( .D(N271), .CP(clk), .CD(rst), .Q(regA[2]) );
  CFD2QX2 \regA_reg[3]  ( .D(N272), .CP(clk), .CD(rst), .Q(regA[3]) );
  CFD2QX2 \regA_reg[5]  ( .D(N274), .CP(clk), .CD(rst), .Q(regA[5]) );
  CFD2QX2 \regA_reg[6]  ( .D(N275), .CP(clk), .CD(rst), .Q(regA[6]) );
  CFD2QX2 \regA_reg[7]  ( .D(N276), .CP(clk), .CD(rst), .Q(regA[7]) );
  CFD2QX2 \regA_reg[9]  ( .D(N278), .CP(clk), .CD(rst), .Q(regA[9]) );
  CFD2QX2 \regA_reg[10]  ( .D(N279), .CP(clk), .CD(rst), .Q(regA[10]) );
  CFD2QX2 \regA_reg[11]  ( .D(N280), .CP(clk), .CD(rst), .Q(regA[11]) );
  CFD2QX2 \regA_reg[16]  ( .D(N285), .CP(clk), .CD(rst), .Q(regA[16]) );
  CFD2QX2 \regA_reg[19]  ( .D(N288), .CP(clk), .CD(rst), .Q(regA[19]) );
  CFD2QX2 \regA_reg[22]  ( .D(N291), .CP(clk), .CD(rst), .Q(regA[22]) );
  CFD2QX2 \regA_reg[23]  ( .D(N292), .CP(clk), .CD(rst), .Q(regA[23]) );
  CFD2QX2 \regA_reg[28]  ( .D(N297), .CP(clk), .CD(rst), .Q(regA[28]) );
  nios_2_DW01_add_8 add_152_4 ( .A({regA[31:30], n2029, regA[28], n2071, n2015, 
        n2036, n2058, regA[23:21], n1379, regA[19], n2126, n2025, regA[16:15], 
        n1494, regA[13], n1475, regA[11:9], n2059, regA[7:2], n2108, n1388}), 
        .B({regB[31:24], n2021, regB[22:18], n2051, n2106, regB[15:14], n2026, 
        regB[12], n2033, regB[10:6], n2049, n2110, n1685, n2047, regB[1:0]}), 
        .CI(1'b0), .SUM({N168, N167, N166, N165, N164, N163, N162, N161, N160, 
        N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, 
        N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137}) );
  nios_2_DW01_add_6 add_152 ( .A({regA[31:30], n2029, regA[28], n2071, n2015, 
        n2036, n2058, regA[23:21], n1379, regA[19], n2125, n2024, regA[16:15], 
        n1494, regA[13], n1475, regA[11:9], n2059, regA[7:2], n2108, n1387}), 
        .B({immi_val[31:11], n2118, immi_val[9:5], n2061, immi_val[3:0]}), 
        .CI(1'b0), .SUM({N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, 
        N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, 
        N70, N69, N68, N67, N66, N65, N64}) );
  nios_2_DW01_add_10 add_152_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, prog_count_ex[7:2], N129, N128}), .B({
        immi_val[31:11], n2118, immi_val[9:5], n2061, immi_val[3:0]}), .CI(
        1'b0), .SUM({N127, N126, N125, N124, N123, N122, N121, N120, N119, 
        N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, 
        N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96}) );
  nios_2_DW01_cmp6_2 r69 ( .A({regB[31:24], n2020, regB[22:18], n2051, n2106, 
        regB[15:14], n2026, regB[12], n2033, regB[10:6], n2049, n2110, n1685, 
        n2047, regB[1:0]}), .B({regA[31:30], n2029, regA[28], n2071, n2015, 
        n2036, n2057, regA[23:21], n1379, regA[19], n2125, n2024, regA[16:15], 
        n1494, regA[13], n1475, regA[11:9], n2059, regA[7:2], n2108, n1387}), 
        .TC(1'b0), .GT(N30), .EQ(N32), .NE(N31) );
  nios_2_DW01_sub_3 sub_152 ( .A({regA[31:30], n2029, regA[28], n2071, n2016, 
        n2037, n2058, regA[23:21], n1380, regA[19], n2126, n2025, regA[16:15], 
        n1495, regA[13], n1476, regA[11:9], n2059, regA[7:2], n2109, n1388}), 
        .B({\twos_comp[31] , \twos_comp[30] , \twos_comp[29] , \twos_comp[28] , 
        \twos_comp[27] , \twos_comp[26] , \twos_comp[25] , \twos_comp[24] , 
        \twos_comp[23] , \twos_comp[22] , \twos_comp[21] , \twos_comp[20] , 
        \twos_comp[19] , \twos_comp[18] , \twos_comp[17] , \twos_comp[16] , 
        \twos_comp[15] , \twos_comp[14] , \twos_comp[13] , \twos_comp[12] , 
        \twos_comp[11] , \twos_comp[10] , \twos_comp[9] , \twos_comp[8] , 
        \twos_comp[7] , \twos_comp[6] , \twos_comp[5] , \twos_comp[4] , 
        \twos_comp[3] , \twos_comp[2] , \twos_comp[1] , \twos_comp[0] }), .CI(
        1'b0), .DIFF({N200, N199, N198, N197, N196, N195, N194, N193, N192, 
        N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, 
        N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169}) );
  nios_2_DW01_inc_3 add_150 ( .A({n5246, \dp_cluster_0/N33 , 
        \dp_cluster_0/N34 , \dp_cluster_0/N35 , \dp_cluster_0/N36 , 
        \dp_cluster_0/N37 , \dp_cluster_0/N38 , \dp_cluster_0/N39 , 
        \dp_cluster_0/N40 , \dp_cluster_0/N41 , \dp_cluster_0/N42 , 
        \dp_cluster_0/N43 , \dp_cluster_0/N44 , \dp_cluster_0/N45 , 
        \dp_cluster_0/N46 , \dp_cluster_0/N47 , \dp_cluster_0/N48 , 
        \dp_cluster_0/N49 , \dp_cluster_0/N50 , \dp_cluster_0/N51 , 
        \dp_cluster_0/N52 , n2119, \dp_cluster_0/N54 , \dp_cluster_0/N55 , 
        \dp_cluster_0/N56 , \dp_cluster_0/N57 , \dp_cluster_0/N58 , n2062, 
        \dp_cluster_0/N60 , \dp_cluster_0/N61 , \dp_cluster_0/N62 , 
        \dp_cluster_0/N63 }), .SUM({\twos_comp[31] , \twos_comp[30] , 
        \twos_comp[29] , \twos_comp[28] , \twos_comp[27] , \twos_comp[26] , 
        \twos_comp[25] , \twos_comp[24] , \twos_comp[23] , \twos_comp[22] , 
        \twos_comp[21] , \twos_comp[20] , \twos_comp[19] , \twos_comp[18] , 
        \twos_comp[17] , \twos_comp[16] , \twos_comp[15] , \twos_comp[14] , 
        \twos_comp[13] , \twos_comp[12] , \twos_comp[11] , \twos_comp[10] , 
        \twos_comp[9] , \twos_comp[8] , \twos_comp[7] , \twos_comp[6] , 
        \twos_comp[5] , \twos_comp[4] , \twos_comp[3] , \twos_comp[2] , 
        \twos_comp[1] , \twos_comp[0] }) );
  CFD2QXL \reg_mem_reg[2][29]  ( .D(n1282), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][29] ) );
  CFD2QXL \reg_mem_reg[0][8]  ( .D(n1367), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][8] ) );
  CFD2QXL \reg_mem_reg[1][8]  ( .D(n1335), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][8] ) );
  CFD2QXL \reg_mem_reg[8][25]  ( .D(n1094), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][25] ) );
  CFD2QXL \reg_mem_reg[4][29]  ( .D(n1218), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][29] ) );
  CFD2QXL \opcode_ex_reg[0]  ( .D(net87782), .CP(clk), .CD(rst), .Q(
        opcode_ex[0]) );
  CFD2QXL \opcode_ex_reg[1]  ( .D(net88155), .CP(clk), .CD(rst), .Q(
        opcode_ex[1]) );
  CFD1QXL \reg_mem_reg[21][15]  ( .D(n688), .CP(clk), .Q(\reg_mem[21][15] ) );
  CFD1QXL \reg_mem_reg[21][21]  ( .D(n682), .CP(clk), .Q(\reg_mem[21][21] ) );
  CFD1QXL \reg_mem_reg[13][15]  ( .D(n944), .CP(clk), .Q(\reg_mem[13][15] ) );
  CFD1QXL \reg_mem_reg[13][21]  ( .D(n938), .CP(clk), .Q(\reg_mem[13][21] ) );
  CFD1QXL \reg_mem_reg[28][15]  ( .D(n464), .CP(clk), .Q(\reg_mem[28][15] ) );
  CFD1QXL \reg_mem_reg[28][21]  ( .D(n458), .CP(clk), .Q(\reg_mem[28][21] ) );
  CFD1QXL \reg_mem_reg[20][31]  ( .D(n704), .CP(clk), .Q(\reg_mem[20][31] ) );
  CFD1QXL \reg_mem_reg[12][15]  ( .D(n976), .CP(clk), .Q(\reg_mem[12][15] ) );
  CFD1QXL \reg_mem_reg[12][21]  ( .D(n970), .CP(clk), .Q(\reg_mem[12][21] ) );
  CFD1QXL \reg_mem_reg[27][15]  ( .D(n496), .CP(clk), .Q(\reg_mem[27][15] ) );
  CFD1QXL \reg_mem_reg[27][21]  ( .D(n490), .CP(clk), .Q(\reg_mem[27][21] ) );
  CFD1QXL \reg_mem_reg[19][15]  ( .D(n752), .CP(clk), .Q(\reg_mem[19][15] ) );
  CFD1QXL \reg_mem_reg[19][21]  ( .D(n746), .CP(clk), .Q(\reg_mem[19][21] ) );
  CFD1QXL \reg_mem_reg[11][15]  ( .D(n1008), .CP(clk), .Q(\reg_mem[11][15] )
         );
  CFD1QXL \reg_mem_reg[11][21]  ( .D(n1002), .CP(clk), .Q(\reg_mem[11][21] )
         );
  CFD1QXL \reg_mem_reg[26][15]  ( .D(n528), .CP(clk), .Q(\reg_mem[26][15] ) );
  CFD1QXL \reg_mem_reg[26][21]  ( .D(n522), .CP(clk), .Q(\reg_mem[26][21] ) );
  CFD1QXL \reg_mem_reg[10][15]  ( .D(n1040), .CP(clk), .Q(\reg_mem[10][15] )
         );
  CFD1QXL \reg_mem_reg[10][21]  ( .D(n1034), .CP(clk), .Q(\reg_mem[10][21] )
         );
  CFD1QXL \reg_mem_reg[23][15]  ( .D(n624), .CP(clk), .Q(\reg_mem[23][15] ) );
  CFD1QXL \reg_mem_reg[23][21]  ( .D(n618), .CP(clk), .Q(\reg_mem[23][21] ) );
  CFD1QXL \reg_mem_reg[15][15]  ( .D(n880), .CP(clk), .Q(\reg_mem[15][15] ) );
  CFD1QXL \reg_mem_reg[15][21]  ( .D(n874), .CP(clk), .Q(\reg_mem[15][21] ) );
  CFD1QXL \reg_mem_reg[22][31]  ( .D(n640), .CP(clk), .Q(\reg_mem[22][31] ) );
  CFD1QXL \reg_mem_reg[14][15]  ( .D(n912), .CP(clk), .Q(\reg_mem[14][15] ) );
  CFD1QXL \reg_mem_reg[14][21]  ( .D(n906), .CP(clk), .Q(\reg_mem[14][21] ) );
  CFD1QXL \reg_mem_reg[25][15]  ( .D(n560), .CP(clk), .Q(\reg_mem[25][15] ) );
  CFD1QXL \reg_mem_reg[25][21]  ( .D(n554), .CP(clk), .Q(\reg_mem[25][21] ) );
  CFD1QXL \reg_mem_reg[17][15]  ( .D(n816), .CP(clk), .Q(\reg_mem[17][15] ) );
  CFD1QXL \reg_mem_reg[17][21]  ( .D(n810), .CP(clk), .Q(\reg_mem[17][21] ) );
  CFD1QXL \reg_mem_reg[24][15]  ( .D(n592), .CP(clk), .Q(\reg_mem[24][15] ) );
  CFD1QXL \reg_mem_reg[24][21]  ( .D(n586), .CP(clk), .Q(\reg_mem[24][21] ) );
  CFD1QXL \reg_mem_reg[21][0]  ( .D(n703), .CP(clk), .Q(\reg_mem[21][0] ) );
  CFD1QXL \reg_mem_reg[21][1]  ( .D(n702), .CP(clk), .Q(\reg_mem[21][1] ) );
  CFD1QXL \reg_mem_reg[21][2]  ( .D(n701), .CP(clk), .Q(\reg_mem[21][2] ) );
  CFD1QXL \reg_mem_reg[21][3]  ( .D(n700), .CP(clk), .Q(\reg_mem[21][3] ) );
  CFD1QXL \reg_mem_reg[21][4]  ( .D(n699), .CP(clk), .Q(\reg_mem[21][4] ) );
  CFD1QXL \reg_mem_reg[21][5]  ( .D(n698), .CP(clk), .Q(\reg_mem[21][5] ) );
  CFD1QXL \reg_mem_reg[21][6]  ( .D(n697), .CP(clk), .Q(\reg_mem[21][6] ) );
  CFD1QXL \reg_mem_reg[21][7]  ( .D(n696), .CP(clk), .Q(\reg_mem[21][7] ) );
  CFD1QXL \reg_mem_reg[21][8]  ( .D(n695), .CP(clk), .Q(\reg_mem[21][8] ) );
  CFD1QXL \reg_mem_reg[21][9]  ( .D(n694), .CP(clk), .Q(\reg_mem[21][9] ) );
  CFD1QXL \reg_mem_reg[21][10]  ( .D(n693), .CP(clk), .Q(\reg_mem[21][10] ) );
  CFD1QXL \reg_mem_reg[21][11]  ( .D(n692), .CP(clk), .Q(\reg_mem[21][11] ) );
  CFD1QXL \reg_mem_reg[21][12]  ( .D(n691), .CP(clk), .Q(\reg_mem[21][12] ) );
  CFD1QXL \reg_mem_reg[21][13]  ( .D(n690), .CP(clk), .Q(\reg_mem[21][13] ) );
  CFD1QXL \reg_mem_reg[21][18]  ( .D(n685), .CP(clk), .Q(\reg_mem[21][18] ) );
  CFD1QXL \reg_mem_reg[21][24]  ( .D(n679), .CP(clk), .Q(\reg_mem[21][24] ) );
  CFD1QXL \reg_mem_reg[21][27]  ( .D(n676), .CP(clk), .Q(\reg_mem[21][27] ) );
  CFD1QXL \reg_mem_reg[21][28]  ( .D(n675), .CP(clk), .Q(\reg_mem[21][28] ) );
  CFD1QXL \reg_mem_reg[21][29]  ( .D(n674), .CP(clk), .Q(\reg_mem[21][29] ) );
  CFD1QXL \reg_mem_reg[21][30]  ( .D(n673), .CP(clk), .Q(\reg_mem[21][30] ) );
  CFD1QXL \reg_mem_reg[21][31]  ( .D(n672), .CP(clk), .Q(\reg_mem[21][31] ) );
  CFD1QXL \reg_mem_reg[13][0]  ( .D(n959), .CP(clk), .Q(\reg_mem[13][0] ) );
  CFD1QXL \reg_mem_reg[13][1]  ( .D(n958), .CP(clk), .Q(\reg_mem[13][1] ) );
  CFD1QXL \reg_mem_reg[13][2]  ( .D(n957), .CP(clk), .Q(\reg_mem[13][2] ) );
  CFD1QXL \reg_mem_reg[13][3]  ( .D(n956), .CP(clk), .Q(\reg_mem[13][3] ) );
  CFD1QXL \reg_mem_reg[13][4]  ( .D(n955), .CP(clk), .Q(\reg_mem[13][4] ) );
  CFD1QXL \reg_mem_reg[13][5]  ( .D(n954), .CP(clk), .Q(\reg_mem[13][5] ) );
  CFD1QXL \reg_mem_reg[13][6]  ( .D(n953), .CP(clk), .Q(\reg_mem[13][6] ) );
  CFD1QXL \reg_mem_reg[13][7]  ( .D(n952), .CP(clk), .Q(\reg_mem[13][7] ) );
  CFD1QXL \reg_mem_reg[13][8]  ( .D(n951), .CP(clk), .Q(\reg_mem[13][8] ) );
  CFD1QXL \reg_mem_reg[13][9]  ( .D(n950), .CP(clk), .Q(\reg_mem[13][9] ) );
  CFD1QXL \reg_mem_reg[13][10]  ( .D(n949), .CP(clk), .Q(\reg_mem[13][10] ) );
  CFD1QXL \reg_mem_reg[13][11]  ( .D(n948), .CP(clk), .Q(\reg_mem[13][11] ) );
  CFD1QXL \reg_mem_reg[13][12]  ( .D(n947), .CP(clk), .Q(\reg_mem[13][12] ) );
  CFD1QXL \reg_mem_reg[13][13]  ( .D(n946), .CP(clk), .Q(\reg_mem[13][13] ) );
  CFD1QXL \reg_mem_reg[13][14]  ( .D(n945), .CP(clk), .Q(\reg_mem[13][14] ) );
  CFD1QXL \reg_mem_reg[13][16]  ( .D(n943), .CP(clk), .Q(\reg_mem[13][16] ) );
  CFD1QXL \reg_mem_reg[13][17]  ( .D(n942), .CP(clk), .Q(\reg_mem[13][17] ) );
  CFD1QXL \reg_mem_reg[13][19]  ( .D(n940), .CP(clk), .Q(\reg_mem[13][19] ) );
  CFD1QXL \reg_mem_reg[28][12]  ( .D(n467), .CP(clk), .Q(\reg_mem[28][12] ) );
  CFD1QXL \reg_mem_reg[28][13]  ( .D(n466), .CP(clk), .Q(\reg_mem[28][13] ) );
  CFD1QXL \reg_mem_reg[28][14]  ( .D(n465), .CP(clk), .Q(\reg_mem[28][14] ) );
  CFD1QXL \reg_mem_reg[28][16]  ( .D(n463), .CP(clk), .Q(\reg_mem[28][16] ) );
  CFD1QXL \reg_mem_reg[28][17]  ( .D(n462), .CP(clk), .Q(\reg_mem[28][17] ) );
  CFD1QXL \reg_mem_reg[28][18]  ( .D(n461), .CP(clk), .Q(\reg_mem[28][18] ) );
  CFD1QXL \reg_mem_reg[28][19]  ( .D(n460), .CP(clk), .Q(\reg_mem[28][19] ) );
  CFD1QXL \reg_mem_reg[28][24]  ( .D(n455), .CP(clk), .Q(\reg_mem[28][24] ) );
  CFD1QXL \reg_mem_reg[28][27]  ( .D(n452), .CP(clk), .Q(\reg_mem[28][27] ) );
  CFD1QXL \reg_mem_reg[28][28]  ( .D(n451), .CP(clk), .Q(\reg_mem[28][28] ) );
  CFD1QXL \reg_mem_reg[28][29]  ( .D(n450), .CP(clk), .Q(\reg_mem[28][29] ) );
  CFD1QXL \reg_mem_reg[28][30]  ( .D(n449), .CP(clk), .Q(\reg_mem[28][30] ) );
  CFD1QXL \reg_mem_reg[28][31]  ( .D(n448), .CP(clk), .Q(\reg_mem[28][31] ) );
  CFD1QXL \reg_mem_reg[20][12]  ( .D(n723), .CP(clk), .Q(\reg_mem[20][12] ) );
  CFD1QXL \reg_mem_reg[20][13]  ( .D(n722), .CP(clk), .Q(\reg_mem[20][13] ) );
  CFD1QXL \reg_mem_reg[20][15]  ( .D(n720), .CP(clk), .Q(\reg_mem[20][15] ) );
  CFD1QXL \reg_mem_reg[20][18]  ( .D(n717), .CP(clk), .Q(\reg_mem[20][18] ) );
  CFD1QXL \reg_mem_reg[20][21]  ( .D(n714), .CP(clk), .Q(\reg_mem[20][21] ) );
  CFD1QXL \reg_mem_reg[20][24]  ( .D(n711), .CP(clk), .Q(\reg_mem[20][24] ) );
  CFD1QXL \reg_mem_reg[20][27]  ( .D(n708), .CP(clk), .Q(\reg_mem[20][27] ) );
  CFD1QXL \reg_mem_reg[20][28]  ( .D(n707), .CP(clk), .Q(\reg_mem[20][28] ) );
  CFD1QXL \reg_mem_reg[20][30]  ( .D(n705), .CP(clk), .Q(\reg_mem[20][30] ) );
  CFD1QXL \reg_mem_reg[12][1]  ( .D(n990), .CP(clk), .Q(\reg_mem[12][1] ) );
  CFD1QXL \reg_mem_reg[12][11]  ( .D(n980), .CP(clk), .Q(\reg_mem[12][11] ) );
  CFD1QXL \reg_mem_reg[12][12]  ( .D(n979), .CP(clk), .Q(\reg_mem[12][12] ) );
  CFD1QXL \reg_mem_reg[12][13]  ( .D(n978), .CP(clk), .Q(\reg_mem[12][13] ) );
  CFD1QXL \reg_mem_reg[12][14]  ( .D(n977), .CP(clk), .Q(\reg_mem[12][14] ) );
  CFD1QXL \reg_mem_reg[12][16]  ( .D(n975), .CP(clk), .Q(\reg_mem[12][16] ) );
  CFD1QXL \reg_mem_reg[12][17]  ( .D(n974), .CP(clk), .Q(\reg_mem[12][17] ) );
  CFD1QXL \reg_mem_reg[12][19]  ( .D(n972), .CP(clk), .Q(\reg_mem[12][19] ) );
  CFD1QXL \reg_mem_reg[27][0]  ( .D(n511), .CP(clk), .Q(\reg_mem[27][0] ) );
  CFD1QXL \reg_mem_reg[27][1]  ( .D(n510), .CP(clk), .Q(\reg_mem[27][1] ) );
  CFD1QXL \reg_mem_reg[27][2]  ( .D(n509), .CP(clk), .Q(\reg_mem[27][2] ) );
  CFD1QXL \reg_mem_reg[27][3]  ( .D(n508), .CP(clk), .Q(\reg_mem[27][3] ) );
  CFD1QXL \reg_mem_reg[27][4]  ( .D(n507), .CP(clk), .Q(\reg_mem[27][4] ) );
  CFD1QXL \reg_mem_reg[27][5]  ( .D(n506), .CP(clk), .Q(\reg_mem[27][5] ) );
  CFD1QXL \reg_mem_reg[27][6]  ( .D(n505), .CP(clk), .Q(\reg_mem[27][6] ) );
  CFD1QXL \reg_mem_reg[27][7]  ( .D(n504), .CP(clk), .Q(\reg_mem[27][7] ) );
  CFD1QXL \reg_mem_reg[27][8]  ( .D(n503), .CP(clk), .Q(\reg_mem[27][8] ) );
  CFD1QXL \reg_mem_reg[27][9]  ( .D(n502), .CP(clk), .Q(\reg_mem[27][9] ) );
  CFD1QXL \reg_mem_reg[27][10]  ( .D(n501), .CP(clk), .Q(\reg_mem[27][10] ) );
  CFD1QXL \reg_mem_reg[27][11]  ( .D(n500), .CP(clk), .Q(\reg_mem[27][11] ) );
  CFD1QXL \reg_mem_reg[27][14]  ( .D(n497), .CP(clk), .Q(\reg_mem[27][14] ) );
  CFD1QXL \reg_mem_reg[27][16]  ( .D(n495), .CP(clk), .Q(\reg_mem[27][16] ) );
  CFD1QXL \reg_mem_reg[27][17]  ( .D(n494), .CP(clk), .Q(\reg_mem[27][17] ) );
  CFD1QXL \reg_mem_reg[27][18]  ( .D(n493), .CP(clk), .Q(\reg_mem[27][18] ) );
  CFD1QXL \reg_mem_reg[27][19]  ( .D(n492), .CP(clk), .Q(\reg_mem[27][19] ) );
  CFD1QXL \reg_mem_reg[27][24]  ( .D(n487), .CP(clk), .Q(\reg_mem[27][24] ) );
  CFD1QXL \reg_mem_reg[27][27]  ( .D(n484), .CP(clk), .Q(\reg_mem[27][27] ) );
  CFD1QXL \reg_mem_reg[27][28]  ( .D(n483), .CP(clk), .Q(\reg_mem[27][28] ) );
  CFD1QXL \reg_mem_reg[27][29]  ( .D(n482), .CP(clk), .Q(\reg_mem[27][29] ) );
  CFD1QXL \reg_mem_reg[27][30]  ( .D(n481), .CP(clk), .Q(\reg_mem[27][30] ) );
  CFD1QXL \reg_mem_reg[27][31]  ( .D(n480), .CP(clk), .Q(\reg_mem[27][31] ) );
  CFD1QXL \reg_mem_reg[19][0]  ( .D(n767), .CP(clk), .Q(\reg_mem[19][0] ) );
  CFD1QXL \reg_mem_reg[19][1]  ( .D(n766), .CP(clk), .Q(\reg_mem[19][1] ) );
  CFD1QXL \reg_mem_reg[19][2]  ( .D(n765), .CP(clk), .Q(\reg_mem[19][2] ) );
  CFD1QXL \reg_mem_reg[19][3]  ( .D(n764), .CP(clk), .Q(\reg_mem[19][3] ) );
  CFD1QXL \reg_mem_reg[19][4]  ( .D(n763), .CP(clk), .Q(\reg_mem[19][4] ) );
  CFD1QXL \reg_mem_reg[19][5]  ( .D(n762), .CP(clk), .Q(\reg_mem[19][5] ) );
  CFD1QXL \reg_mem_reg[19][6]  ( .D(n761), .CP(clk), .Q(\reg_mem[19][6] ) );
  CFD1QXL \reg_mem_reg[19][7]  ( .D(n760), .CP(clk), .Q(\reg_mem[19][7] ) );
  CFD1QXL \reg_mem_reg[19][8]  ( .D(n759), .CP(clk), .Q(\reg_mem[19][8] ) );
  CFD1QXL \reg_mem_reg[19][9]  ( .D(n758), .CP(clk), .Q(\reg_mem[19][9] ) );
  CFD1QXL \reg_mem_reg[19][10]  ( .D(n757), .CP(clk), .Q(\reg_mem[19][10] ) );
  CFD1QXL \reg_mem_reg[19][11]  ( .D(n756), .CP(clk), .Q(\reg_mem[19][11] ) );
  CFD1QXL \reg_mem_reg[19][18]  ( .D(n749), .CP(clk), .Q(\reg_mem[19][18] ) );
  CFD1QXL \reg_mem_reg[19][24]  ( .D(n743), .CP(clk), .Q(\reg_mem[19][24] ) );
  CFD1QXL \reg_mem_reg[19][27]  ( .D(n740), .CP(clk), .Q(\reg_mem[19][27] ) );
  CFD1QXL \reg_mem_reg[19][28]  ( .D(n739), .CP(clk), .Q(\reg_mem[19][28] ) );
  CFD1QXL \reg_mem_reg[19][29]  ( .D(n738), .CP(clk), .Q(\reg_mem[19][29] ) );
  CFD1QXL \reg_mem_reg[19][30]  ( .D(n737), .CP(clk), .Q(\reg_mem[19][30] ) );
  CFD1QXL \reg_mem_reg[19][31]  ( .D(n736), .CP(clk), .Q(\reg_mem[19][31] ) );
  CFD1QXL \reg_mem_reg[11][0]  ( .D(n1023), .CP(clk), .Q(\reg_mem[11][0] ) );
  CFD1QXL \reg_mem_reg[11][2]  ( .D(n1021), .CP(clk), .Q(\reg_mem[11][2] ) );
  CFD1QXL \reg_mem_reg[11][3]  ( .D(n1020), .CP(clk), .Q(\reg_mem[11][3] ) );
  CFD1QXL \reg_mem_reg[11][4]  ( .D(n1019), .CP(clk), .Q(\reg_mem[11][4] ) );
  CFD1QXL \reg_mem_reg[11][5]  ( .D(n1018), .CP(clk), .Q(\reg_mem[11][5] ) );
  CFD1QXL \reg_mem_reg[11][6]  ( .D(n1017), .CP(clk), .Q(\reg_mem[11][6] ) );
  CFD1QXL \reg_mem_reg[11][7]  ( .D(n1016), .CP(clk), .Q(\reg_mem[11][7] ) );
  CFD1QXL \reg_mem_reg[11][8]  ( .D(n1015), .CP(clk), .Q(\reg_mem[11][8] ) );
  CFD1QXL \reg_mem_reg[11][9]  ( .D(n1014), .CP(clk), .Q(\reg_mem[11][9] ) );
  CFD1QXL \reg_mem_reg[11][10]  ( .D(n1013), .CP(clk), .Q(\reg_mem[11][10] )
         );
  CFD1QXL \reg_mem_reg[11][13]  ( .D(n1010), .CP(clk), .Q(\reg_mem[11][13] )
         );
  CFD1QXL \reg_mem_reg[11][14]  ( .D(n1009), .CP(clk), .Q(\reg_mem[11][14] )
         );
  CFD1QXL \reg_mem_reg[11][16]  ( .D(n1007), .CP(clk), .Q(\reg_mem[11][16] )
         );
  CFD1QXL \reg_mem_reg[11][17]  ( .D(n1006), .CP(clk), .Q(\reg_mem[11][17] )
         );
  CFD1QXL \reg_mem_reg[11][19]  ( .D(n1004), .CP(clk), .Q(\reg_mem[11][19] )
         );
  CFD1QXL \reg_mem_reg[26][14]  ( .D(n529), .CP(clk), .Q(\reg_mem[26][14] ) );
  CFD1QXL \reg_mem_reg[26][16]  ( .D(n527), .CP(clk), .Q(\reg_mem[26][16] ) );
  CFD1QXL \reg_mem_reg[26][17]  ( .D(n526), .CP(clk), .Q(\reg_mem[26][17] ) );
  CFD1QXL \reg_mem_reg[26][18]  ( .D(n525), .CP(clk), .Q(\reg_mem[26][18] ) );
  CFD1QXL \reg_mem_reg[26][19]  ( .D(n524), .CP(clk), .Q(\reg_mem[26][19] ) );
  CFD1QXL \reg_mem_reg[26][24]  ( .D(n519), .CP(clk), .Q(\reg_mem[26][24] ) );
  CFD1QXL \reg_mem_reg[26][27]  ( .D(n516), .CP(clk), .Q(\reg_mem[26][27] ) );
  CFD1QXL \reg_mem_reg[26][28]  ( .D(n515), .CP(clk), .Q(\reg_mem[26][28] ) );
  CFD1QXL \reg_mem_reg[26][29]  ( .D(n514), .CP(clk), .Q(\reg_mem[26][29] ) );
  CFD1QXL \reg_mem_reg[26][30]  ( .D(n513), .CP(clk), .Q(\reg_mem[26][30] ) );
  CFD1QXL \reg_mem_reg[26][31]  ( .D(n512), .CP(clk), .Q(\reg_mem[26][31] ) );
  CFD1QXL \reg_mem_reg[18][15]  ( .D(n784), .CP(clk), .Q(\reg_mem[18][15] ) );
  CFD1QXL \reg_mem_reg[18][18]  ( .D(n781), .CP(clk), .Q(\reg_mem[18][18] ) );
  CFD1QXL \reg_mem_reg[18][21]  ( .D(n778), .CP(clk), .Q(\reg_mem[18][21] ) );
  CFD1QXL \reg_mem_reg[18][24]  ( .D(n775), .CP(clk), .Q(\reg_mem[18][24] ) );
  CFD1QXL \reg_mem_reg[18][27]  ( .D(n772), .CP(clk), .Q(\reg_mem[18][27] ) );
  CFD1QXL \reg_mem_reg[18][28]  ( .D(n771), .CP(clk), .Q(\reg_mem[18][28] ) );
  CFD1QXL \reg_mem_reg[18][30]  ( .D(n769), .CP(clk), .Q(\reg_mem[18][30] ) );
  CFD1QXL \reg_mem_reg[10][13]  ( .D(n1042), .CP(clk), .Q(\reg_mem[10][13] )
         );
  CFD1QXL \reg_mem_reg[10][14]  ( .D(n1041), .CP(clk), .Q(\reg_mem[10][14] )
         );
  CFD1QXL \reg_mem_reg[10][16]  ( .D(n1039), .CP(clk), .Q(\reg_mem[10][16] )
         );
  CFD1QXL \reg_mem_reg[10][17]  ( .D(n1038), .CP(clk), .Q(\reg_mem[10][17] )
         );
  CFD1QXL \reg_mem_reg[10][19]  ( .D(n1036), .CP(clk), .Q(\reg_mem[10][19] )
         );
  CFD1QXL \reg_mem_reg[23][0]  ( .D(n639), .CP(clk), .Q(\reg_mem[23][0] ) );
  CFD1QXL \reg_mem_reg[23][1]  ( .D(n638), .CP(clk), .Q(\reg_mem[23][1] ) );
  CFD1QXL \reg_mem_reg[23][2]  ( .D(n637), .CP(clk), .Q(\reg_mem[23][2] ) );
  CFD1QXL \reg_mem_reg[23][3]  ( .D(n636), .CP(clk), .Q(\reg_mem[23][3] ) );
  CFD1QXL \reg_mem_reg[23][4]  ( .D(n635), .CP(clk), .Q(\reg_mem[23][4] ) );
  CFD1QXL \reg_mem_reg[23][5]  ( .D(n634), .CP(clk), .Q(\reg_mem[23][5] ) );
  CFD1QXL \reg_mem_reg[23][6]  ( .D(n633), .CP(clk), .Q(\reg_mem[23][6] ) );
  CFD1QXL \reg_mem_reg[23][7]  ( .D(n632), .CP(clk), .Q(\reg_mem[23][7] ) );
  CFD1QXL \reg_mem_reg[23][8]  ( .D(n631), .CP(clk), .Q(\reg_mem[23][8] ) );
  CFD1QXL \reg_mem_reg[23][9]  ( .D(n630), .CP(clk), .Q(\reg_mem[23][9] ) );
  CFD1QXL \reg_mem_reg[23][10]  ( .D(n629), .CP(clk), .Q(\reg_mem[23][10] ) );
  CFD1QXL \reg_mem_reg[23][11]  ( .D(n628), .CP(clk), .Q(\reg_mem[23][11] ) );
  CFD1QXL \reg_mem_reg[23][12]  ( .D(n627), .CP(clk), .Q(\reg_mem[23][12] ) );
  CFD1QXL \reg_mem_reg[23][13]  ( .D(n626), .CP(clk), .Q(\reg_mem[23][13] ) );
  CFD1QXL \reg_mem_reg[23][18]  ( .D(n621), .CP(clk), .Q(\reg_mem[23][18] ) );
  CFD1QXL \reg_mem_reg[23][24]  ( .D(n615), .CP(clk), .Q(\reg_mem[23][24] ) );
  CFD1QXL \reg_mem_reg[23][27]  ( .D(n612), .CP(clk), .Q(\reg_mem[23][27] ) );
  CFD1QXL \reg_mem_reg[23][28]  ( .D(n611), .CP(clk), .Q(\reg_mem[23][28] ) );
  CFD1QXL \reg_mem_reg[23][29]  ( .D(n610), .CP(clk), .Q(\reg_mem[23][29] ) );
  CFD1QXL \reg_mem_reg[23][30]  ( .D(n609), .CP(clk), .Q(\reg_mem[23][30] ) );
  CFD1QXL \reg_mem_reg[23][31]  ( .D(n608), .CP(clk), .Q(\reg_mem[23][31] ) );
  CFD1QXL \reg_mem_reg[15][0]  ( .D(n895), .CP(clk), .Q(\reg_mem[15][0] ) );
  CFD1QXL \reg_mem_reg[15][2]  ( .D(n893), .CP(clk), .Q(\reg_mem[15][2] ) );
  CFD1QXL \reg_mem_reg[15][3]  ( .D(n892), .CP(clk), .Q(\reg_mem[15][3] ) );
  CFD1QXL \reg_mem_reg[15][4]  ( .D(n891), .CP(clk), .Q(\reg_mem[15][4] ) );
  CFD1QXL \reg_mem_reg[15][5]  ( .D(n890), .CP(clk), .Q(\reg_mem[15][5] ) );
  CFD1QXL \reg_mem_reg[15][6]  ( .D(n889), .CP(clk), .Q(\reg_mem[15][6] ) );
  CFD1QXL \reg_mem_reg[15][7]  ( .D(n888), .CP(clk), .Q(\reg_mem[15][7] ) );
  CFD1QXL \reg_mem_reg[15][8]  ( .D(n887), .CP(clk), .Q(\reg_mem[15][8] ) );
  CFD1QXL \reg_mem_reg[15][9]  ( .D(n886), .CP(clk), .Q(\reg_mem[15][9] ) );
  CFD1QXL \reg_mem_reg[15][10]  ( .D(n885), .CP(clk), .Q(\reg_mem[15][10] ) );
  CFD1QXL \reg_mem_reg[15][11]  ( .D(n884), .CP(clk), .Q(\reg_mem[15][11] ) );
  CFD1QXL \reg_mem_reg[15][12]  ( .D(n883), .CP(clk), .Q(\reg_mem[15][12] ) );
  CFD1QXL \reg_mem_reg[15][13]  ( .D(n882), .CP(clk), .Q(\reg_mem[15][13] ) );
  CFD1QXL \reg_mem_reg[15][14]  ( .D(n881), .CP(clk), .Q(\reg_mem[15][14] ) );
  CFD1QXL \reg_mem_reg[15][16]  ( .D(n879), .CP(clk), .Q(\reg_mem[15][16] ) );
  CFD1QXL \reg_mem_reg[15][17]  ( .D(n878), .CP(clk), .Q(\reg_mem[15][17] ) );
  CFD1QXL \reg_mem_reg[15][19]  ( .D(n876), .CP(clk), .Q(\reg_mem[15][19] ) );
  CFD1QXL \reg_mem_reg[22][12]  ( .D(n659), .CP(clk), .Q(\reg_mem[22][12] ) );
  CFD1QXL \reg_mem_reg[22][13]  ( .D(n658), .CP(clk), .Q(\reg_mem[22][13] ) );
  CFD1QXL \reg_mem_reg[22][15]  ( .D(n656), .CP(clk), .Q(\reg_mem[22][15] ) );
  CFD1QXL \reg_mem_reg[22][18]  ( .D(n653), .CP(clk), .Q(\reg_mem[22][18] ) );
  CFD1QXL \reg_mem_reg[22][21]  ( .D(n650), .CP(clk), .Q(\reg_mem[22][21] ) );
  CFD1QXL \reg_mem_reg[22][24]  ( .D(n647), .CP(clk), .Q(\reg_mem[22][24] ) );
  CFD1QXL \reg_mem_reg[22][27]  ( .D(n644), .CP(clk), .Q(\reg_mem[22][27] ) );
  CFD1QXL \reg_mem_reg[22][28]  ( .D(n643), .CP(clk), .Q(\reg_mem[22][28] ) );
  CFD1QXL \reg_mem_reg[22][29]  ( .D(n642), .CP(clk), .Q(\reg_mem[22][29] ) );
  CFD1QXL \reg_mem_reg[22][30]  ( .D(n641), .CP(clk), .Q(\reg_mem[22][30] ) );
  CFD1QXL \reg_mem_reg[14][1]  ( .D(n926), .CP(clk), .Q(\reg_mem[14][1] ) );
  CFD1QXL \reg_mem_reg[14][11]  ( .D(n916), .CP(clk), .Q(\reg_mem[14][11] ) );
  CFD1QXL \reg_mem_reg[14][12]  ( .D(n915), .CP(clk), .Q(\reg_mem[14][12] ) );
  CFD1QXL \reg_mem_reg[14][13]  ( .D(n914), .CP(clk), .Q(\reg_mem[14][13] ) );
  CFD1QXL \reg_mem_reg[14][14]  ( .D(n913), .CP(clk), .Q(\reg_mem[14][14] ) );
  CFD1QXL \reg_mem_reg[14][16]  ( .D(n911), .CP(clk), .Q(\reg_mem[14][16] ) );
  CFD1QXL \reg_mem_reg[14][17]  ( .D(n910), .CP(clk), .Q(\reg_mem[14][17] ) );
  CFD1QXL \reg_mem_reg[14][19]  ( .D(n908), .CP(clk), .Q(\reg_mem[14][19] ) );
  CFD1QXL \reg_mem_reg[25][0]  ( .D(n575), .CP(clk), .Q(\reg_mem[25][0] ) );
  CFD1QXL \reg_mem_reg[25][1]  ( .D(n574), .CP(clk), .Q(\reg_mem[25][1] ) );
  CFD1QXL \reg_mem_reg[25][2]  ( .D(n573), .CP(clk), .Q(\reg_mem[25][2] ) );
  CFD1QXL \reg_mem_reg[25][3]  ( .D(n572), .CP(clk), .Q(\reg_mem[25][3] ) );
  CFD1QXL \reg_mem_reg[25][4]  ( .D(n571), .CP(clk), .Q(\reg_mem[25][4] ) );
  CFD1QXL \reg_mem_reg[25][5]  ( .D(n570), .CP(clk), .Q(\reg_mem[25][5] ) );
  CFD1QXL \reg_mem_reg[25][6]  ( .D(n569), .CP(clk), .Q(\reg_mem[25][6] ) );
  CFD1QXL \reg_mem_reg[25][7]  ( .D(n568), .CP(clk), .Q(\reg_mem[25][7] ) );
  CFD1QXL \reg_mem_reg[25][8]  ( .D(n567), .CP(clk), .Q(\reg_mem[25][8] ) );
  CFD1QXL \reg_mem_reg[25][9]  ( .D(n566), .CP(clk), .Q(\reg_mem[25][9] ) );
  CFD1QXL \reg_mem_reg[25][10]  ( .D(n565), .CP(clk), .Q(\reg_mem[25][10] ) );
  CFD1QXL \reg_mem_reg[25][11]  ( .D(n564), .CP(clk), .Q(\reg_mem[25][11] ) );
  CFD1QXL \reg_mem_reg[25][14]  ( .D(n561), .CP(clk), .Q(\reg_mem[25][14] ) );
  CFD1QXL \reg_mem_reg[25][16]  ( .D(n559), .CP(clk), .Q(\reg_mem[25][16] ) );
  CFD1QXL \reg_mem_reg[25][17]  ( .D(n558), .CP(clk), .Q(\reg_mem[25][17] ) );
  CFD1QXL \reg_mem_reg[25][18]  ( .D(n557), .CP(clk), .Q(\reg_mem[25][18] ) );
  CFD1QXL \reg_mem_reg[25][19]  ( .D(n556), .CP(clk), .Q(\reg_mem[25][19] ) );
  CFD1QXL \reg_mem_reg[25][24]  ( .D(n551), .CP(clk), .Q(\reg_mem[25][24] ) );
  CFD1QXL \reg_mem_reg[25][27]  ( .D(n548), .CP(clk), .Q(\reg_mem[25][27] ) );
  CFD1QXL \reg_mem_reg[25][28]  ( .D(n547), .CP(clk), .Q(\reg_mem[25][28] ) );
  CFD1QXL \reg_mem_reg[25][29]  ( .D(n546), .CP(clk), .Q(\reg_mem[25][29] ) );
  CFD1QXL \reg_mem_reg[25][30]  ( .D(n545), .CP(clk), .Q(\reg_mem[25][30] ) );
  CFD1QXL \reg_mem_reg[25][31]  ( .D(n544), .CP(clk), .Q(\reg_mem[25][31] ) );
  CFD1QXL \reg_mem_reg[17][0]  ( .D(n831), .CP(clk), .Q(\reg_mem[17][0] ) );
  CFD1QXL \reg_mem_reg[17][1]  ( .D(n830), .CP(clk), .Q(\reg_mem[17][1] ) );
  CFD1QXL \reg_mem_reg[17][2]  ( .D(n829), .CP(clk), .Q(\reg_mem[17][2] ) );
  CFD1QXL \reg_mem_reg[17][3]  ( .D(n828), .CP(clk), .Q(\reg_mem[17][3] ) );
  CFD1QXL \reg_mem_reg[17][4]  ( .D(n827), .CP(clk), .Q(\reg_mem[17][4] ) );
  CFD1QXL \reg_mem_reg[17][5]  ( .D(n826), .CP(clk), .Q(\reg_mem[17][5] ) );
  CFD1QXL \reg_mem_reg[17][6]  ( .D(n825), .CP(clk), .Q(\reg_mem[17][6] ) );
  CFD1QXL \reg_mem_reg[17][7]  ( .D(n824), .CP(clk), .Q(\reg_mem[17][7] ) );
  CFD1QXL \reg_mem_reg[17][8]  ( .D(n823), .CP(clk), .Q(\reg_mem[17][8] ) );
  CFD1QXL \reg_mem_reg[17][9]  ( .D(n822), .CP(clk), .Q(\reg_mem[17][9] ) );
  CFD1QXL \reg_mem_reg[17][10]  ( .D(n821), .CP(clk), .Q(\reg_mem[17][10] ) );
  CFD1QXL \reg_mem_reg[17][11]  ( .D(n820), .CP(clk), .Q(\reg_mem[17][11] ) );
  CFD1QXL \reg_mem_reg[17][18]  ( .D(n813), .CP(clk), .Q(\reg_mem[17][18] ) );
  CFD1QXL \reg_mem_reg[17][24]  ( .D(n807), .CP(clk), .Q(\reg_mem[17][24] ) );
  CFD1QXL \reg_mem_reg[17][27]  ( .D(n804), .CP(clk), .Q(\reg_mem[17][27] ) );
  CFD1QXL \reg_mem_reg[17][28]  ( .D(n803), .CP(clk), .Q(\reg_mem[17][28] ) );
  CFD1QXL \reg_mem_reg[17][30]  ( .D(n801), .CP(clk), .Q(\reg_mem[17][30] ) );
  CFD1QXL \reg_mem_reg[17][31]  ( .D(n800), .CP(clk), .Q(\reg_mem[17][31] ) );
  CFD1QXL \reg_mem_reg[24][14]  ( .D(n593), .CP(clk), .Q(\reg_mem[24][14] ) );
  CFD1QXL \reg_mem_reg[24][16]  ( .D(n591), .CP(clk), .Q(\reg_mem[24][16] ) );
  CFD1QXL \reg_mem_reg[24][17]  ( .D(n590), .CP(clk), .Q(\reg_mem[24][17] ) );
  CFD1QXL \reg_mem_reg[24][18]  ( .D(n589), .CP(clk), .Q(\reg_mem[24][18] ) );
  CFD1QXL \reg_mem_reg[24][19]  ( .D(n588), .CP(clk), .Q(\reg_mem[24][19] ) );
  CFD1QXL \reg_mem_reg[24][24]  ( .D(n583), .CP(clk), .Q(\reg_mem[24][24] ) );
  CFD1QXL \reg_mem_reg[24][27]  ( .D(n580), .CP(clk), .Q(\reg_mem[24][27] ) );
  CFD1QXL \reg_mem_reg[24][28]  ( .D(n579), .CP(clk), .Q(\reg_mem[24][28] ) );
  CFD1QXL \reg_mem_reg[24][29]  ( .D(n578), .CP(clk), .Q(\reg_mem[24][29] ) );
  CFD1QXL \reg_mem_reg[24][30]  ( .D(n577), .CP(clk), .Q(\reg_mem[24][30] ) );
  CFD1QXL \reg_mem_reg[24][31]  ( .D(n576), .CP(clk), .Q(\reg_mem[24][31] ) );
  CFD1QXL \reg_mem_reg[16][15]  ( .D(n848), .CP(clk), .Q(\reg_mem[16][15] ) );
  CFD1QXL \reg_mem_reg[16][18]  ( .D(n845), .CP(clk), .Q(\reg_mem[16][18] ) );
  CFD1QXL \reg_mem_reg[16][21]  ( .D(n842), .CP(clk), .Q(\reg_mem[16][21] ) );
  CFD1QXL \reg_mem_reg[16][24]  ( .D(n839), .CP(clk), .Q(\reg_mem[16][24] ) );
  CFD1QXL \reg_mem_reg[16][27]  ( .D(n836), .CP(clk), .Q(\reg_mem[16][27] ) );
  CFD1QXL \reg_mem_reg[16][28]  ( .D(n835), .CP(clk), .Q(\reg_mem[16][28] ) );
  CFD1QXL \reg_mem_reg[16][29]  ( .D(n834), .CP(clk), .Q(\reg_mem[16][29] ) );
  CFD1QXL \reg_mem_reg[16][30]  ( .D(n833), .CP(clk), .Q(\reg_mem[16][30] ) );
  CFD1QXL \reg_mem_reg[21][14]  ( .D(n689), .CP(clk), .Q(\reg_mem[21][14] ) );
  CFD1QXL \reg_mem_reg[21][16]  ( .D(n687), .CP(clk), .Q(\reg_mem[21][16] ) );
  CFD1QXL \reg_mem_reg[21][17]  ( .D(n686), .CP(clk), .Q(\reg_mem[21][17] ) );
  CFD1QXL \reg_mem_reg[21][19]  ( .D(n684), .CP(clk), .Q(\reg_mem[21][19] ) );
  CFD1QXL \reg_mem_reg[13][18]  ( .D(n941), .CP(clk), .Q(\reg_mem[13][18] ) );
  CFD1QXL \reg_mem_reg[13][24]  ( .D(n935), .CP(clk), .Q(\reg_mem[13][24] ) );
  CFD1QXL \reg_mem_reg[13][27]  ( .D(n932), .CP(clk), .Q(\reg_mem[13][27] ) );
  CFD1QXL \reg_mem_reg[13][28]  ( .D(n931), .CP(clk), .Q(\reg_mem[13][28] ) );
  CFD1QXL \reg_mem_reg[13][29]  ( .D(n930), .CP(clk), .Q(\reg_mem[13][29] ) );
  CFD1QXL \reg_mem_reg[13][30]  ( .D(n929), .CP(clk), .Q(\reg_mem[13][30] ) );
  CFD1QXL \reg_mem_reg[13][31]  ( .D(n928), .CP(clk), .Q(\reg_mem[13][31] ) );
  CFD1QXL \reg_mem_reg[28][0]  ( .D(n479), .CP(clk), .Q(\reg_mem[28][0] ) );
  CFD1QXL \reg_mem_reg[28][1]  ( .D(n478), .CP(clk), .Q(\reg_mem[28][1] ) );
  CFD1QXL \reg_mem_reg[28][2]  ( .D(n477), .CP(clk), .Q(\reg_mem[28][2] ) );
  CFD1QXL \reg_mem_reg[28][3]  ( .D(n476), .CP(clk), .Q(\reg_mem[28][3] ) );
  CFD1QXL \reg_mem_reg[28][4]  ( .D(n475), .CP(clk), .Q(\reg_mem[28][4] ) );
  CFD1QXL \reg_mem_reg[28][5]  ( .D(n474), .CP(clk), .Q(\reg_mem[28][5] ) );
  CFD1QXL \reg_mem_reg[28][6]  ( .D(n473), .CP(clk), .Q(\reg_mem[28][6] ) );
  CFD1QXL \reg_mem_reg[28][7]  ( .D(n472), .CP(clk), .Q(\reg_mem[28][7] ) );
  CFD1QXL \reg_mem_reg[28][8]  ( .D(n471), .CP(clk), .Q(\reg_mem[28][8] ) );
  CFD1QXL \reg_mem_reg[28][9]  ( .D(n470), .CP(clk), .Q(\reg_mem[28][9] ) );
  CFD1QXL \reg_mem_reg[28][10]  ( .D(n469), .CP(clk), .Q(\reg_mem[28][10] ) );
  CFD1QXL \reg_mem_reg[28][11]  ( .D(n468), .CP(clk), .Q(\reg_mem[28][11] ) );
  CFD1QXL \reg_mem_reg[20][0]  ( .D(n735), .CP(clk), .Q(\reg_mem[20][0] ) );
  CFD1QXL \reg_mem_reg[20][1]  ( .D(n734), .CP(clk), .Q(\reg_mem[20][1] ) );
  CFD1QXL \reg_mem_reg[20][2]  ( .D(n733), .CP(clk), .Q(\reg_mem[20][2] ) );
  CFD1QXL \reg_mem_reg[20][3]  ( .D(n732), .CP(clk), .Q(\reg_mem[20][3] ) );
  CFD1QXL \reg_mem_reg[20][4]  ( .D(n731), .CP(clk), .Q(\reg_mem[20][4] ) );
  CFD1QXL \reg_mem_reg[20][5]  ( .D(n730), .CP(clk), .Q(\reg_mem[20][5] ) );
  CFD1QXL \reg_mem_reg[20][6]  ( .D(n729), .CP(clk), .Q(\reg_mem[20][6] ) );
  CFD1QXL \reg_mem_reg[20][7]  ( .D(n728), .CP(clk), .Q(\reg_mem[20][7] ) );
  CFD1QXL \reg_mem_reg[20][8]  ( .D(n727), .CP(clk), .Q(\reg_mem[20][8] ) );
  CFD1QXL \reg_mem_reg[20][9]  ( .D(n726), .CP(clk), .Q(\reg_mem[20][9] ) );
  CFD1QXL \reg_mem_reg[20][10]  ( .D(n725), .CP(clk), .Q(\reg_mem[20][10] ) );
  CFD1QXL \reg_mem_reg[20][11]  ( .D(n724), .CP(clk), .Q(\reg_mem[20][11] ) );
  CFD1QXL \reg_mem_reg[20][14]  ( .D(n721), .CP(clk), .Q(\reg_mem[20][14] ) );
  CFD1QXL \reg_mem_reg[20][16]  ( .D(n719), .CP(clk), .Q(\reg_mem[20][16] ) );
  CFD1QXL \reg_mem_reg[20][17]  ( .D(n718), .CP(clk), .Q(\reg_mem[20][17] ) );
  CFD1QXL \reg_mem_reg[20][19]  ( .D(n716), .CP(clk), .Q(\reg_mem[20][19] ) );
  CFD1QXL \reg_mem_reg[12][0]  ( .D(n991), .CP(clk), .Q(\reg_mem[12][0] ) );
  CFD1QXL \reg_mem_reg[12][2]  ( .D(n989), .CP(clk), .Q(\reg_mem[12][2] ) );
  CFD1QXL \reg_mem_reg[12][3]  ( .D(n988), .CP(clk), .Q(\reg_mem[12][3] ) );
  CFD1QXL \reg_mem_reg[12][4]  ( .D(n987), .CP(clk), .Q(\reg_mem[12][4] ) );
  CFD1QXL \reg_mem_reg[12][5]  ( .D(n986), .CP(clk), .Q(\reg_mem[12][5] ) );
  CFD1QXL \reg_mem_reg[12][6]  ( .D(n985), .CP(clk), .Q(\reg_mem[12][6] ) );
  CFD1QXL \reg_mem_reg[12][7]  ( .D(n984), .CP(clk), .Q(\reg_mem[12][7] ) );
  CFD1QXL \reg_mem_reg[12][8]  ( .D(n983), .CP(clk), .Q(\reg_mem[12][8] ) );
  CFD1QXL \reg_mem_reg[12][9]  ( .D(n982), .CP(clk), .Q(\reg_mem[12][9] ) );
  CFD1QXL \reg_mem_reg[12][10]  ( .D(n981), .CP(clk), .Q(\reg_mem[12][10] ) );
  CFD1QXL \reg_mem_reg[12][18]  ( .D(n973), .CP(clk), .Q(\reg_mem[12][18] ) );
  CFD1QXL \reg_mem_reg[12][24]  ( .D(n967), .CP(clk), .Q(\reg_mem[12][24] ) );
  CFD1QXL \reg_mem_reg[12][27]  ( .D(n964), .CP(clk), .Q(\reg_mem[12][27] ) );
  CFD1QXL \reg_mem_reg[12][28]  ( .D(n963), .CP(clk), .Q(\reg_mem[12][28] ) );
  CFD1QXL \reg_mem_reg[12][29]  ( .D(n962), .CP(clk), .Q(\reg_mem[12][29] ) );
  CFD1QXL \reg_mem_reg[12][30]  ( .D(n961), .CP(clk), .Q(\reg_mem[12][30] ) );
  CFD1QXL \reg_mem_reg[12][31]  ( .D(n960), .CP(clk), .Q(\reg_mem[12][31] ) );
  CFD1QXL \reg_mem_reg[27][12]  ( .D(n499), .CP(clk), .Q(\reg_mem[27][12] ) );
  CFD1QXL \reg_mem_reg[27][13]  ( .D(n498), .CP(clk), .Q(\reg_mem[27][13] ) );
  CFD1QXL \reg_mem_reg[19][12]  ( .D(n755), .CP(clk), .Q(\reg_mem[19][12] ) );
  CFD1QXL \reg_mem_reg[19][13]  ( .D(n754), .CP(clk), .Q(\reg_mem[19][13] ) );
  CFD1QXL \reg_mem_reg[19][14]  ( .D(n753), .CP(clk), .Q(\reg_mem[19][14] ) );
  CFD1QXL \reg_mem_reg[19][16]  ( .D(n751), .CP(clk), .Q(\reg_mem[19][16] ) );
  CFD1QXL \reg_mem_reg[19][17]  ( .D(n750), .CP(clk), .Q(\reg_mem[19][17] ) );
  CFD1QXL \reg_mem_reg[19][19]  ( .D(n748), .CP(clk), .Q(\reg_mem[19][19] ) );
  CFD1QXL \reg_mem_reg[11][11]  ( .D(n1012), .CP(clk), .Q(\reg_mem[11][11] )
         );
  CFD1QXL \reg_mem_reg[11][12]  ( .D(n1011), .CP(clk), .Q(\reg_mem[11][12] )
         );
  CFD1QXL \reg_mem_reg[11][18]  ( .D(n1005), .CP(clk), .Q(\reg_mem[11][18] )
         );
  CFD1QXL \reg_mem_reg[11][24]  ( .D(n999), .CP(clk), .Q(\reg_mem[11][24] ) );
  CFD1QXL \reg_mem_reg[11][27]  ( .D(n996), .CP(clk), .Q(\reg_mem[11][27] ) );
  CFD1QXL \reg_mem_reg[11][28]  ( .D(n995), .CP(clk), .Q(\reg_mem[11][28] ) );
  CFD1QXL \reg_mem_reg[11][29]  ( .D(n994), .CP(clk), .Q(\reg_mem[11][29] ) );
  CFD1QXL \reg_mem_reg[11][30]  ( .D(n993), .CP(clk), .Q(\reg_mem[11][30] ) );
  CFD1QXL \reg_mem_reg[11][31]  ( .D(n992), .CP(clk), .Q(\reg_mem[11][31] ) );
  CFD1QXL \reg_mem_reg[26][0]  ( .D(n543), .CP(clk), .Q(\reg_mem[26][0] ) );
  CFD1QXL \reg_mem_reg[26][1]  ( .D(n542), .CP(clk), .Q(\reg_mem[26][1] ) );
  CFD1QXL \reg_mem_reg[26][2]  ( .D(n541), .CP(clk), .Q(\reg_mem[26][2] ) );
  CFD1QXL \reg_mem_reg[26][3]  ( .D(n540), .CP(clk), .Q(\reg_mem[26][3] ) );
  CFD1QXL \reg_mem_reg[26][4]  ( .D(n539), .CP(clk), .Q(\reg_mem[26][4] ) );
  CFD1QXL \reg_mem_reg[26][5]  ( .D(n538), .CP(clk), .Q(\reg_mem[26][5] ) );
  CFD1QXL \reg_mem_reg[26][6]  ( .D(n537), .CP(clk), .Q(\reg_mem[26][6] ) );
  CFD1QXL \reg_mem_reg[26][7]  ( .D(n536), .CP(clk), .Q(\reg_mem[26][7] ) );
  CFD1QXL \reg_mem_reg[26][8]  ( .D(n535), .CP(clk), .Q(\reg_mem[26][8] ) );
  CFD1QXL \reg_mem_reg[26][9]  ( .D(n534), .CP(clk), .Q(\reg_mem[26][9] ) );
  CFD1QXL \reg_mem_reg[26][10]  ( .D(n533), .CP(clk), .Q(\reg_mem[26][10] ) );
  CFD1QXL \reg_mem_reg[26][11]  ( .D(n532), .CP(clk), .Q(\reg_mem[26][11] ) );
  CFD1QXL \reg_mem_reg[26][12]  ( .D(n531), .CP(clk), .Q(\reg_mem[26][12] ) );
  CFD1QXL \reg_mem_reg[26][13]  ( .D(n530), .CP(clk), .Q(\reg_mem[26][13] ) );
  CFD1QXL \reg_mem_reg[18][0]  ( .D(n799), .CP(clk), .Q(\reg_mem[18][0] ) );
  CFD1QXL \reg_mem_reg[18][1]  ( .D(n798), .CP(clk), .Q(\reg_mem[18][1] ) );
  CFD1QXL \reg_mem_reg[18][2]  ( .D(n797), .CP(clk), .Q(\reg_mem[18][2] ) );
  CFD1QXL \reg_mem_reg[18][3]  ( .D(n796), .CP(clk), .Q(\reg_mem[18][3] ) );
  CFD1QXL \reg_mem_reg[18][4]  ( .D(n795), .CP(clk), .Q(\reg_mem[18][4] ) );
  CFD1QXL \reg_mem_reg[18][5]  ( .D(n794), .CP(clk), .Q(\reg_mem[18][5] ) );
  CFD1QXL \reg_mem_reg[18][6]  ( .D(n793), .CP(clk), .Q(\reg_mem[18][6] ) );
  CFD1QXL \reg_mem_reg[18][7]  ( .D(n792), .CP(clk), .Q(\reg_mem[18][7] ) );
  CFD1QXL \reg_mem_reg[18][8]  ( .D(n791), .CP(clk), .Q(\reg_mem[18][8] ) );
  CFD1QXL \reg_mem_reg[18][9]  ( .D(n790), .CP(clk), .Q(\reg_mem[18][9] ) );
  CFD1QXL \reg_mem_reg[18][10]  ( .D(n789), .CP(clk), .Q(\reg_mem[18][10] ) );
  CFD1QXL \reg_mem_reg[18][11]  ( .D(n788), .CP(clk), .Q(\reg_mem[18][11] ) );
  CFD1QXL \reg_mem_reg[18][12]  ( .D(n787), .CP(clk), .Q(\reg_mem[18][12] ) );
  CFD1QXL \reg_mem_reg[18][13]  ( .D(n786), .CP(clk), .Q(\reg_mem[18][13] ) );
  CFD1QXL \reg_mem_reg[18][14]  ( .D(n785), .CP(clk), .Q(\reg_mem[18][14] ) );
  CFD1QXL \reg_mem_reg[18][16]  ( .D(n783), .CP(clk), .Q(\reg_mem[18][16] ) );
  CFD1QXL \reg_mem_reg[18][17]  ( .D(n782), .CP(clk), .Q(\reg_mem[18][17] ) );
  CFD1QXL \reg_mem_reg[18][19]  ( .D(n780), .CP(clk), .Q(\reg_mem[18][19] ) );
  CFD1QXL \reg_mem_reg[10][0]  ( .D(n1055), .CP(clk), .Q(\reg_mem[10][0] ) );
  CFD1QXL \reg_mem_reg[10][1]  ( .D(n1054), .CP(clk), .Q(\reg_mem[10][1] ) );
  CFD1QXL \reg_mem_reg[10][2]  ( .D(n1053), .CP(clk), .Q(\reg_mem[10][2] ) );
  CFD1QXL \reg_mem_reg[10][3]  ( .D(n1052), .CP(clk), .Q(\reg_mem[10][3] ) );
  CFD1QXL \reg_mem_reg[10][4]  ( .D(n1051), .CP(clk), .Q(\reg_mem[10][4] ) );
  CFD1QXL \reg_mem_reg[10][5]  ( .D(n1050), .CP(clk), .Q(\reg_mem[10][5] ) );
  CFD1QXL \reg_mem_reg[10][6]  ( .D(n1049), .CP(clk), .Q(\reg_mem[10][6] ) );
  CFD1QXL \reg_mem_reg[10][7]  ( .D(n1048), .CP(clk), .Q(\reg_mem[10][7] ) );
  CFD1QXL \reg_mem_reg[10][8]  ( .D(n1047), .CP(clk), .Q(\reg_mem[10][8] ) );
  CFD1QXL \reg_mem_reg[10][9]  ( .D(n1046), .CP(clk), .Q(\reg_mem[10][9] ) );
  CFD1QXL \reg_mem_reg[10][10]  ( .D(n1045), .CP(clk), .Q(\reg_mem[10][10] )
         );
  CFD1QXL \reg_mem_reg[10][11]  ( .D(n1044), .CP(clk), .Q(\reg_mem[10][11] )
         );
  CFD1QXL \reg_mem_reg[10][12]  ( .D(n1043), .CP(clk), .Q(\reg_mem[10][12] )
         );
  CFD1QXL \reg_mem_reg[10][18]  ( .D(n1037), .CP(clk), .Q(\reg_mem[10][18] )
         );
  CFD1QXL \reg_mem_reg[10][24]  ( .D(n1031), .CP(clk), .Q(\reg_mem[10][24] )
         );
  CFD1QXL \reg_mem_reg[10][27]  ( .D(n1028), .CP(clk), .Q(\reg_mem[10][27] )
         );
  CFD1QXL \reg_mem_reg[10][28]  ( .D(n1027), .CP(clk), .Q(\reg_mem[10][28] )
         );
  CFD1QXL \reg_mem_reg[10][29]  ( .D(n1026), .CP(clk), .Q(\reg_mem[10][29] )
         );
  CFD1QXL \reg_mem_reg[10][30]  ( .D(n1025), .CP(clk), .Q(\reg_mem[10][30] )
         );
  CFD1QXL \reg_mem_reg[10][31]  ( .D(n1024), .CP(clk), .Q(\reg_mem[10][31] )
         );
  CFD1QXL \reg_mem_reg[23][14]  ( .D(n625), .CP(clk), .Q(\reg_mem[23][14] ) );
  CFD1QXL \reg_mem_reg[23][16]  ( .D(n623), .CP(clk), .Q(\reg_mem[23][16] ) );
  CFD1QXL \reg_mem_reg[23][17]  ( .D(n622), .CP(clk), .Q(\reg_mem[23][17] ) );
  CFD1QXL \reg_mem_reg[23][19]  ( .D(n620), .CP(clk), .Q(\reg_mem[23][19] ) );
  CFD1QXL \reg_mem_reg[15][18]  ( .D(n877), .CP(clk), .Q(\reg_mem[15][18] ) );
  CFD1QXL \reg_mem_reg[15][24]  ( .D(n871), .CP(clk), .Q(\reg_mem[15][24] ) );
  CFD1QXL \reg_mem_reg[15][27]  ( .D(n868), .CP(clk), .Q(\reg_mem[15][27] ) );
  CFD1QXL \reg_mem_reg[15][28]  ( .D(n867), .CP(clk), .Q(\reg_mem[15][28] ) );
  CFD1QXL \reg_mem_reg[15][29]  ( .D(n866), .CP(clk), .Q(\reg_mem[15][29] ) );
  CFD1QXL \reg_mem_reg[15][30]  ( .D(n865), .CP(clk), .Q(\reg_mem[15][30] ) );
  CFD1QXL \reg_mem_reg[15][31]  ( .D(n864), .CP(clk), .Q(\reg_mem[15][31] ) );
  CFD1QXL \reg_mem_reg[22][0]  ( .D(n671), .CP(clk), .Q(\reg_mem[22][0] ) );
  CFD1QXL \reg_mem_reg[22][1]  ( .D(n670), .CP(clk), .Q(\reg_mem[22][1] ) );
  CFD1QXL \reg_mem_reg[22][2]  ( .D(n669), .CP(clk), .Q(\reg_mem[22][2] ) );
  CFD1QXL \reg_mem_reg[22][3]  ( .D(n668), .CP(clk), .Q(\reg_mem[22][3] ) );
  CFD1QXL \reg_mem_reg[22][4]  ( .D(n667), .CP(clk), .Q(\reg_mem[22][4] ) );
  CFD1QXL \reg_mem_reg[22][5]  ( .D(n666), .CP(clk), .Q(\reg_mem[22][5] ) );
  CFD1QXL \reg_mem_reg[22][6]  ( .D(n665), .CP(clk), .Q(\reg_mem[22][6] ) );
  CFD1QXL \reg_mem_reg[22][7]  ( .D(n664), .CP(clk), .Q(\reg_mem[22][7] ) );
  CFD1QXL \reg_mem_reg[22][8]  ( .D(n663), .CP(clk), .Q(\reg_mem[22][8] ) );
  CFD1QXL \reg_mem_reg[22][9]  ( .D(n662), .CP(clk), .Q(\reg_mem[22][9] ) );
  CFD1QXL \reg_mem_reg[22][10]  ( .D(n661), .CP(clk), .Q(\reg_mem[22][10] ) );
  CFD1QXL \reg_mem_reg[22][11]  ( .D(n660), .CP(clk), .Q(\reg_mem[22][11] ) );
  CFD1QXL \reg_mem_reg[22][14]  ( .D(n657), .CP(clk), .Q(\reg_mem[22][14] ) );
  CFD1QXL \reg_mem_reg[22][16]  ( .D(n655), .CP(clk), .Q(\reg_mem[22][16] ) );
  CFD1QXL \reg_mem_reg[22][17]  ( .D(n654), .CP(clk), .Q(\reg_mem[22][17] ) );
  CFD1QXL \reg_mem_reg[22][19]  ( .D(n652), .CP(clk), .Q(\reg_mem[22][19] ) );
  CFD1QXL \reg_mem_reg[14][0]  ( .D(n927), .CP(clk), .Q(\reg_mem[14][0] ) );
  CFD1QXL \reg_mem_reg[14][2]  ( .D(n925), .CP(clk), .Q(\reg_mem[14][2] ) );
  CFD1QXL \reg_mem_reg[14][3]  ( .D(n924), .CP(clk), .Q(\reg_mem[14][3] ) );
  CFD1QXL \reg_mem_reg[14][4]  ( .D(n923), .CP(clk), .Q(\reg_mem[14][4] ) );
  CFD1QXL \reg_mem_reg[14][5]  ( .D(n922), .CP(clk), .Q(\reg_mem[14][5] ) );
  CFD1QXL \reg_mem_reg[14][6]  ( .D(n921), .CP(clk), .Q(\reg_mem[14][6] ) );
  CFD1QXL \reg_mem_reg[14][7]  ( .D(n920), .CP(clk), .Q(\reg_mem[14][7] ) );
  CFD1QXL \reg_mem_reg[14][8]  ( .D(n919), .CP(clk), .Q(\reg_mem[14][8] ) );
  CFD1QXL \reg_mem_reg[14][9]  ( .D(n918), .CP(clk), .Q(\reg_mem[14][9] ) );
  CFD1QXL \reg_mem_reg[14][10]  ( .D(n917), .CP(clk), .Q(\reg_mem[14][10] ) );
  CFD1QXL \reg_mem_reg[14][18]  ( .D(n909), .CP(clk), .Q(\reg_mem[14][18] ) );
  CFD1QXL \reg_mem_reg[14][24]  ( .D(n903), .CP(clk), .Q(\reg_mem[14][24] ) );
  CFD1QXL \reg_mem_reg[14][27]  ( .D(n900), .CP(clk), .Q(\reg_mem[14][27] ) );
  CFD1QXL \reg_mem_reg[14][28]  ( .D(n899), .CP(clk), .Q(\reg_mem[14][28] ) );
  CFD1QXL \reg_mem_reg[14][29]  ( .D(n898), .CP(clk), .Q(\reg_mem[14][29] ) );
  CFD1QXL \reg_mem_reg[14][30]  ( .D(n897), .CP(clk), .Q(\reg_mem[14][30] ) );
  CFD1QXL \reg_mem_reg[14][31]  ( .D(n896), .CP(clk), .Q(\reg_mem[14][31] ) );
  CFD1QXL \reg_mem_reg[25][12]  ( .D(n563), .CP(clk), .Q(\reg_mem[25][12] ) );
  CFD1QXL \reg_mem_reg[25][13]  ( .D(n562), .CP(clk), .Q(\reg_mem[25][13] ) );
  CFD1QXL \reg_mem_reg[17][12]  ( .D(n819), .CP(clk), .Q(\reg_mem[17][12] ) );
  CFD1QXL \reg_mem_reg[17][13]  ( .D(n818), .CP(clk), .Q(\reg_mem[17][13] ) );
  CFD1QXL \reg_mem_reg[17][14]  ( .D(n817), .CP(clk), .Q(\reg_mem[17][14] ) );
  CFD1QXL \reg_mem_reg[17][16]  ( .D(n815), .CP(clk), .Q(\reg_mem[17][16] ) );
  CFD1QXL \reg_mem_reg[17][17]  ( .D(n814), .CP(clk), .Q(\reg_mem[17][17] ) );
  CFD1QXL \reg_mem_reg[17][19]  ( .D(n812), .CP(clk), .Q(\reg_mem[17][19] ) );
  CFD1QXL \reg_mem_reg[24][0]  ( .D(n607), .CP(clk), .Q(\reg_mem[24][0] ) );
  CFD1QXL \reg_mem_reg[24][1]  ( .D(n606), .CP(clk), .Q(\reg_mem[24][1] ) );
  CFD1QXL \reg_mem_reg[24][2]  ( .D(n605), .CP(clk), .Q(\reg_mem[24][2] ) );
  CFD1QXL \reg_mem_reg[24][3]  ( .D(n604), .CP(clk), .Q(\reg_mem[24][3] ) );
  CFD1QXL \reg_mem_reg[24][4]  ( .D(n603), .CP(clk), .Q(\reg_mem[24][4] ) );
  CFD1QXL \reg_mem_reg[24][5]  ( .D(n602), .CP(clk), .Q(\reg_mem[24][5] ) );
  CFD1QXL \reg_mem_reg[24][6]  ( .D(n601), .CP(clk), .Q(\reg_mem[24][6] ) );
  CFD1QXL \reg_mem_reg[24][7]  ( .D(n600), .CP(clk), .Q(\reg_mem[24][7] ) );
  CFD1QXL \reg_mem_reg[24][8]  ( .D(n599), .CP(clk), .Q(\reg_mem[24][8] ) );
  CFD1QXL \reg_mem_reg[24][9]  ( .D(n598), .CP(clk), .Q(\reg_mem[24][9] ) );
  CFD1QXL \reg_mem_reg[24][10]  ( .D(n597), .CP(clk), .Q(\reg_mem[24][10] ) );
  CFD1QXL \reg_mem_reg[24][11]  ( .D(n596), .CP(clk), .Q(\reg_mem[24][11] ) );
  CFD1QXL \reg_mem_reg[24][12]  ( .D(n595), .CP(clk), .Q(\reg_mem[24][12] ) );
  CFD1QXL \reg_mem_reg[24][13]  ( .D(n594), .CP(clk), .Q(\reg_mem[24][13] ) );
  CFD1QXL \reg_mem_reg[16][0]  ( .D(n863), .CP(clk), .Q(\reg_mem[16][0] ) );
  CFD1QXL \reg_mem_reg[16][1]  ( .D(n862), .CP(clk), .Q(\reg_mem[16][1] ) );
  CFD1QXL \reg_mem_reg[16][2]  ( .D(n861), .CP(clk), .Q(\reg_mem[16][2] ) );
  CFD1QXL \reg_mem_reg[16][3]  ( .D(n860), .CP(clk), .Q(\reg_mem[16][3] ) );
  CFD1QXL \reg_mem_reg[16][4]  ( .D(n859), .CP(clk), .Q(\reg_mem[16][4] ) );
  CFD1QXL \reg_mem_reg[16][5]  ( .D(n858), .CP(clk), .Q(\reg_mem[16][5] ) );
  CFD1QXL \reg_mem_reg[16][6]  ( .D(n857), .CP(clk), .Q(\reg_mem[16][6] ) );
  CFD1QXL \reg_mem_reg[16][7]  ( .D(n856), .CP(clk), .Q(\reg_mem[16][7] ) );
  CFD1QXL \reg_mem_reg[16][8]  ( .D(n855), .CP(clk), .Q(\reg_mem[16][8] ) );
  CFD1QXL \reg_mem_reg[16][9]  ( .D(n854), .CP(clk), .Q(\reg_mem[16][9] ) );
  CFD1QXL \reg_mem_reg[16][10]  ( .D(n853), .CP(clk), .Q(\reg_mem[16][10] ) );
  CFD1QXL \reg_mem_reg[16][11]  ( .D(n852), .CP(clk), .Q(\reg_mem[16][11] ) );
  CFD1QXL \reg_mem_reg[16][12]  ( .D(n851), .CP(clk), .Q(\reg_mem[16][12] ) );
  CFD1QXL \reg_mem_reg[16][13]  ( .D(n850), .CP(clk), .Q(\reg_mem[16][13] ) );
  CFD1QXL \reg_mem_reg[16][14]  ( .D(n849), .CP(clk), .Q(\reg_mem[16][14] ) );
  CFD1QXL \reg_mem_reg[16][16]  ( .D(n847), .CP(clk), .Q(\reg_mem[16][16] ) );
  CFD1QXL \reg_mem_reg[16][17]  ( .D(n846), .CP(clk), .Q(\reg_mem[16][17] ) );
  CFD1QXL \reg_mem_reg[16][19]  ( .D(n844), .CP(clk), .Q(\reg_mem[16][19] ) );
  CFD2QXL i_type_mem_reg ( .D(n1692), .CP(clk), .CD(rst), .Q(i_type_mem) );
  CFD2QXL j_type_mem_reg ( .D(n1694), .CP(clk), .CD(rst), .Q(j_type_mem) );
  CFD2QXL \regB_mem_reg[31]  ( .D(n1696), .CP(clk), .CD(rst), .Q(regB_mem[31])
         );
  CFD2QXL \regB_mem_reg[30]  ( .D(n1461), .CP(clk), .CD(rst), .Q(regB_mem[30])
         );
  CFD2QXL \regB_mem_reg[29]  ( .D(n1701), .CP(clk), .CD(rst), .Q(regB_mem[29])
         );
  CFD2QXL \regB_mem_reg[28]  ( .D(n1702), .CP(clk), .CD(rst), .Q(regB_mem[28])
         );
  CFD2QXL \regB_mem_reg[27]  ( .D(n1705), .CP(clk), .CD(rst), .Q(regB_mem[27])
         );
  CFD2QXL \regB_mem_reg[26]  ( .D(n1708), .CP(clk), .CD(rst), .Q(regB_mem[26])
         );
  CFD2QXL \regB_mem_reg[25]  ( .D(n1711), .CP(clk), .CD(rst), .Q(regB_mem[25])
         );
  CFD2QXL \regB_mem_reg[24]  ( .D(n1714), .CP(clk), .CD(rst), .Q(regB_mem[24])
         );
  CFD2QXL \regB_mem_reg[23]  ( .D(n1717), .CP(clk), .CD(rst), .Q(regB_mem[23])
         );
  CFD2QXL \regB_mem_reg[22]  ( .D(n1718), .CP(clk), .CD(rst), .Q(regB_mem[22])
         );
  CFD2QXL \regB_mem_reg[21]  ( .D(n1721), .CP(clk), .CD(rst), .Q(regB_mem[21])
         );
  CFD2QXL \regB_mem_reg[20]  ( .D(n1724), .CP(clk), .CD(rst), .Q(regB_mem[20])
         );
  CFD2QXL \regB_mem_reg[19]  ( .D(n1727), .CP(clk), .CD(rst), .Q(regB_mem[19])
         );
  CFD2QXL \regB_mem_reg[18]  ( .D(n1462), .CP(clk), .CD(rst), .Q(regB_mem[18])
         );
  CFD2QXL \regB_mem_reg[17]  ( .D(n1730), .CP(clk), .CD(rst), .Q(regB_mem[17])
         );
  CFD2QXL \regB_mem_reg[16]  ( .D(n1732), .CP(clk), .CD(rst), .Q(regB_mem[16])
         );
  CFD2QXL \regB_mem_reg[15]  ( .D(n1734), .CP(clk), .CD(rst), .Q(regB_mem[15])
         );
  CFD2QXL \regB_mem_reg[14]  ( .D(n1465), .CP(clk), .CD(rst), .Q(regB_mem[14])
         );
  CFD2QXL \regB_mem_reg[13]  ( .D(n1739), .CP(clk), .CD(rst), .Q(regB_mem[13])
         );
  CFD2QXL \regB_mem_reg[12]  ( .D(n1742), .CP(clk), .CD(rst), .Q(regB_mem[12])
         );
  CFD2QXL \regB_mem_reg[11]  ( .D(n1745), .CP(clk), .CD(rst), .Q(regB_mem[11])
         );
  CFD2QXL \regB_mem_reg[10]  ( .D(n1747), .CP(clk), .CD(rst), .Q(regB_mem[10])
         );
  CFD2QXL \regB_mem_reg[9]  ( .D(n1750), .CP(clk), .CD(rst), .Q(regB_mem[9])
         );
  CFD2QXL \regB_mem_reg[8]  ( .D(n1753), .CP(clk), .CD(rst), .Q(regB_mem[8])
         );
  CFD2QXL \regB_mem_reg[7]  ( .D(n1756), .CP(clk), .CD(rst), .Q(regB_mem[7])
         );
  CFD2QXL \regB_mem_reg[6]  ( .D(n1759), .CP(clk), .CD(rst), .Q(regB_mem[6])
         );
  CFD2QXL \regB_mem_reg[5]  ( .D(n1762), .CP(clk), .CD(rst), .Q(regB_mem[5])
         );
  CFD2QXL \regB_mem_reg[4]  ( .D(n1763), .CP(clk), .CD(rst), .Q(regB_mem[4])
         );
  CFD2QXL \regB_mem_reg[3]  ( .D(n1765), .CP(clk), .CD(rst), .Q(regB_mem[3])
         );
  CFD2QXL \regB_mem_reg[2]  ( .D(n1768), .CP(clk), .CD(rst), .Q(regB_mem[2])
         );
  CFD2QXL \regB_mem_reg[1]  ( .D(n1771), .CP(clk), .CD(rst), .Q(regB_mem[1])
         );
  CFD2QXL \regB_mem_reg[0]  ( .D(n1772), .CP(clk), .CD(rst), .Q(regB_mem[0])
         );
  CFD2QXL \alu_op_reg[8]  ( .D(alu_op_c[8]), .CP(clk), .CD(rst), .Q(alu_op[8])
         );
  CFD2QXL \alu_op_reg[31]  ( .D(alu_op_c[31]), .CP(clk), .CD(rst), .Q(
        alu_op[31]) );
  CFD2QXL \alu_op_reg[30]  ( .D(alu_op_c[30]), .CP(clk), .CD(rst), .Q(
        alu_op[30]) );
  CFD2QXL \alu_op_reg[1]  ( .D(alu_op_c[1]), .CP(clk), .CD(rst), .Q(alu_op[1])
         );
  CFD2QXL \alu_op_reg[2]  ( .D(alu_op_c[2]), .CP(clk), .CD(rst), .Q(alu_op[2])
         );
  CFD2QXL \alu_op_reg[3]  ( .D(alu_op_c[3]), .CP(clk), .CD(rst), .Q(alu_op[3])
         );
  CFD2QXL \alu_op_reg[4]  ( .D(alu_op_c[4]), .CP(clk), .CD(rst), .Q(alu_op[4])
         );
  CFD2QXL \alu_op_reg[5]  ( .D(alu_op_c[5]), .CP(clk), .CD(rst), .Q(alu_op[5])
         );
  CFD2QXL \alu_op_reg[6]  ( .D(alu_op_c[6]), .CP(clk), .CD(rst), .Q(alu_op[6])
         );
  CFD2QXL \alu_op_reg[7]  ( .D(alu_op_c[7]), .CP(clk), .CD(rst), .Q(alu_op[7])
         );
  CFD2QXL \alu_op_reg[9]  ( .D(alu_op_c[9]), .CP(clk), .CD(rst), .Q(alu_op[9])
         );
  CFD2QXL \alu_op_reg[10]  ( .D(alu_op_c[10]), .CP(clk), .CD(rst), .Q(
        alu_op[10]) );
  CFD2QXL \alu_op_reg[11]  ( .D(alu_op_c[11]), .CP(clk), .CD(rst), .Q(
        alu_op[11]) );
  CFD2QXL \alu_op_reg[12]  ( .D(alu_op_c[12]), .CP(clk), .CD(rst), .Q(
        alu_op[12]) );
  CFD2QXL \alu_op_reg[13]  ( .D(alu_op_c[13]), .CP(clk), .CD(rst), .Q(
        alu_op[13]) );
  CFD2QXL \alu_op_reg[14]  ( .D(alu_op_c[14]), .CP(clk), .CD(rst), .Q(
        alu_op[14]) );
  CFD2QXL \alu_op_reg[15]  ( .D(n5243), .CP(clk), .CD(rst), .Q(alu_op[15]) );
  CFD2QXL \alu_op_reg[16]  ( .D(alu_op_c[16]), .CP(clk), .CD(rst), .Q(
        alu_op[16]) );
  CFD2QXL \alu_op_reg[17]  ( .D(alu_op_c[17]), .CP(clk), .CD(rst), .Q(
        alu_op[17]) );
  CFD2QXL \alu_op_reg[18]  ( .D(alu_op_c[18]), .CP(clk), .CD(rst), .Q(
        alu_op[18]) );
  CFD2QXL \alu_op_reg[19]  ( .D(alu_op_c[19]), .CP(clk), .CD(rst), .Q(
        alu_op[19]) );
  CFD2QXL \alu_op_reg[20]  ( .D(alu_op_c[20]), .CP(clk), .CD(rst), .Q(
        alu_op[20]) );
  CFD2QXL \alu_op_reg[21]  ( .D(n5244), .CP(clk), .CD(rst), .Q(alu_op[21]) );
  CFD2QXL \alu_op_reg[22]  ( .D(n5245), .CP(clk), .CD(rst), .Q(alu_op[22]) );
  CFD2QXL \alu_op_reg[23]  ( .D(alu_op_c[23]), .CP(clk), .CD(rst), .Q(
        alu_op[23]) );
  CFD2QXL \alu_op_reg[24]  ( .D(alu_op_c[24]), .CP(clk), .CD(rst), .Q(
        alu_op[24]) );
  CFD2QXL \alu_op_reg[25]  ( .D(alu_op_c[25]), .CP(clk), .CD(rst), .Q(
        alu_op[25]) );
  CFD2QXL \alu_op_reg[26]  ( .D(alu_op_c[26]), .CP(clk), .CD(rst), .Q(
        alu_op[26]) );
  CFD2QXL \alu_op_reg[27]  ( .D(alu_op_c[27]), .CP(clk), .CD(rst), .Q(
        alu_op[27]) );
  CFD2QXL \alu_op_reg[28]  ( .D(alu_op_c[28]), .CP(clk), .CD(rst), .Q(
        alu_op[28]) );
  CFD2QXL \alu_op_reg[29]  ( .D(alu_op_c[29]), .CP(clk), .CD(rst), .Q(
        alu_op[29]) );
  CFD2QXL \alu_op_reg[0]  ( .D(alu_op_c[0]), .CP(clk), .CD(rst), .Q(alu_op[0])
         );
  CFD2QXL \alu_op_wb_reg[8]  ( .D(n1775), .CP(clk), .CD(rst), .Q(alu_op_wb[8])
         );
  CFD2QXL \alu_op_wb_reg[31]  ( .D(n1777), .CP(clk), .CD(rst), .Q(
        alu_op_wb[31]) );
  CFD2QXL \alu_op_wb_reg[1]  ( .D(n1779), .CP(clk), .CD(rst), .Q(alu_op_wb[1])
         );
  CFD2QXL \alu_op_wb_reg[2]  ( .D(n1781), .CP(clk), .CD(rst), .Q(alu_op_wb[2])
         );
  CFD2QXL \alu_op_wb_reg[3]  ( .D(n1783), .CP(clk), .CD(rst), .Q(alu_op_wb[3])
         );
  CFD2QXL \alu_op_wb_reg[4]  ( .D(n1785), .CP(clk), .CD(rst), .Q(alu_op_wb[4])
         );
  CFD2QXL \alu_op_wb_reg[5]  ( .D(n1787), .CP(clk), .CD(rst), .Q(alu_op_wb[5])
         );
  CFD2QXL \alu_op_wb_reg[6]  ( .D(n1789), .CP(clk), .CD(rst), .Q(alu_op_wb[6])
         );
  CFD2QXL \alu_op_wb_reg[7]  ( .D(n1791), .CP(clk), .CD(rst), .Q(alu_op_wb[7])
         );
  CFD2QXL \alu_op_wb_reg[9]  ( .D(n1793), .CP(clk), .CD(rst), .Q(alu_op_wb[9])
         );
  CFD2QXL \alu_op_wb_reg[10]  ( .D(n1795), .CP(clk), .CD(rst), .Q(
        alu_op_wb[10]) );
  CFD2QXL \alu_op_wb_reg[11]  ( .D(n1797), .CP(clk), .CD(rst), .Q(
        alu_op_wb[11]) );
  CFD2QXL \alu_op_wb_reg[12]  ( .D(n1799), .CP(clk), .CD(rst), .Q(
        alu_op_wb[12]) );
  CFD2QXL \alu_op_wb_reg[0]  ( .D(n1801), .CP(clk), .CD(rst), .Q(alu_op_wb[0])
         );
  CFD2QXL \alu_op_wb_reg[30]  ( .D(n1803), .CP(clk), .CD(rst), .Q(
        alu_op_wb[30]) );
  CFD2QXL \alu_op_wb_reg[13]  ( .D(n1805), .CP(clk), .CD(rst), .Q(
        alu_op_wb[13]) );
  CFD2QXL \alu_op_wb_reg[14]  ( .D(n1807), .CP(clk), .CD(rst), .Q(
        alu_op_wb[14]) );
  CFD2QXL \alu_op_wb_reg[15]  ( .D(n1809), .CP(clk), .CD(rst), .Q(
        alu_op_wb[15]) );
  CFD2QXL \alu_op_wb_reg[16]  ( .D(n1811), .CP(clk), .CD(rst), .Q(
        alu_op_wb[16]) );
  CFD2QXL \alu_op_wb_reg[17]  ( .D(n1813), .CP(clk), .CD(rst), .Q(
        alu_op_wb[17]) );
  CFD2QXL \alu_op_wb_reg[18]  ( .D(n1815), .CP(clk), .CD(rst), .Q(
        alu_op_wb[18]) );
  CFD2QXL \alu_op_wb_reg[19]  ( .D(n1817), .CP(clk), .CD(rst), .Q(
        alu_op_wb[19]) );
  CFD2QXL \alu_op_wb_reg[20]  ( .D(n1819), .CP(clk), .CD(rst), .Q(
        alu_op_wb[20]) );
  CFD2QXL \alu_op_wb_reg[21]  ( .D(n1821), .CP(clk), .CD(rst), .Q(
        alu_op_wb[21]) );
  CFD2QXL \alu_op_wb_reg[22]  ( .D(n1823), .CP(clk), .CD(rst), .Q(
        alu_op_wb[22]) );
  CFD2QXL \alu_op_wb_reg[23]  ( .D(n1825), .CP(clk), .CD(rst), .Q(
        alu_op_wb[23]) );
  CFD2QXL \alu_op_wb_reg[24]  ( .D(n1827), .CP(clk), .CD(rst), .Q(
        alu_op_wb[24]) );
  CFD2QXL \alu_op_wb_reg[25]  ( .D(n1829), .CP(clk), .CD(rst), .Q(
        alu_op_wb[25]) );
  CFD2QXL \alu_op_wb_reg[26]  ( .D(n1831), .CP(clk), .CD(rst), .Q(
        alu_op_wb[26]) );
  CFD2QXL \alu_op_wb_reg[27]  ( .D(n1833), .CP(clk), .CD(rst), .Q(
        alu_op_wb[27]) );
  CFD2QXL \alu_op_wb_reg[28]  ( .D(n1835), .CP(clk), .CD(rst), .Q(
        alu_op_wb[28]) );
  CFD2QXL \alu_op_wb_reg[29]  ( .D(n1837), .CP(clk), .CD(rst), .Q(
        alu_op_wb[29]) );
  CFD2XL \opcode_mem_reg[5]  ( .D(n1839), .CP(clk), .CD(rst), .QN(n98) );
  CFD2QXL \prog_count_reg[7]  ( .D(prog_count_c[7]), .CP(clk), .CD(rst), .Q(
        prog_count_o[7]) );
  CFD2QXL \opcode_mem_reg[2]  ( .D(n1840), .CP(clk), .CD(rst), .Q(
        opcode_mem[2]) );
  CFD2QXL \reg_mem_reg[5][15]  ( .D(n1200), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][15] ) );
  CFD2QXL \reg_mem_reg[5][21]  ( .D(n1194), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][21] ) );
  CFD2QXL \reg_mem_reg[31][15]  ( .D(n368), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][15] ) );
  CFD2QXL \reg_mem_reg[31][21]  ( .D(n362), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][21] ) );
  CFD2QXL \reg_mem_reg[7][15]  ( .D(n1136), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][15] ) );
  CFD2QXL \reg_mem_reg[7][21]  ( .D(n1130), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][21] ) );
  CFD2QXL \reg_mem_reg[9][15]  ( .D(n1072), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][15] ) );
  CFD2QXL \reg_mem_reg[9][21]  ( .D(n1066), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][21] ) );
  CFD2QXL \prog_count_reg[0]  ( .D(prog_count_c[0]), .CP(clk), .CD(rst), .Q(
        N22) );
  CFD2QXL \prog_count_reg[1]  ( .D(prog_count_c[1]), .CP(clk), .CD(rst), .Q(
        N23) );
  CFD2XL \opcode_mem_reg[4]  ( .D(n1841), .CP(clk), .CD(rst), .QN(n99) );
  CFD2XL \opcode_mem_reg[3]  ( .D(n1842), .CP(clk), .CD(rst), .QN(n100) );
  CFD2QXL \reg_mem_reg[29][16]  ( .D(n431), .CP(clk), .CD(rst), .Q(
        \reg_mem[29][16] ) );
  CFD2QXL \reg_mem_reg[29][17]  ( .D(n430), .CP(clk), .CD(rst), .Q(
        \reg_mem[29][17] ) );
  CFD2QXL \reg_mem_reg[29][18]  ( .D(n429), .CP(clk), .CD(rst), .Q(
        \reg_mem[29][18] ) );
  CFD2QXL \reg_mem_reg[29][19]  ( .D(n428), .CP(clk), .CD(rst), .Q(
        \reg_mem[29][19] ) );
  CFD2QXL \reg_mem_reg[29][24]  ( .D(n423), .CP(clk), .CD(rst), .Q(
        \reg_mem[29][24] ) );
  CFD2QXL \reg_mem_reg[29][27]  ( .D(n420), .CP(clk), .CD(rst), .Q(
        \reg_mem[29][27] ) );
  CFD2QXL \reg_mem_reg[29][28]  ( .D(n419), .CP(clk), .CD(rst), .Q(
        \reg_mem[29][28] ) );
  CFD2QXL \reg_mem_reg[29][30]  ( .D(n417), .CP(clk), .CD(rst), .Q(
        \reg_mem[29][30] ) );
  CFD2QXL \reg_mem_reg[5][0]  ( .D(n1215), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][0] ) );
  CFD2QXL \reg_mem_reg[5][1]  ( .D(n1214), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][1] ) );
  CFD2QXL \reg_mem_reg[5][2]  ( .D(n1213), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][2] ) );
  CFD2QXL \reg_mem_reg[5][3]  ( .D(n1212), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][3] ) );
  CFD2QXL \reg_mem_reg[5][4]  ( .D(n1211), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][4] ) );
  CFD2QXL \reg_mem_reg[5][5]  ( .D(n1210), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][5] ) );
  CFD2QXL \reg_mem_reg[5][6]  ( .D(n1209), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][6] ) );
  CFD2QXL \reg_mem_reg[5][7]  ( .D(n1208), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][7] ) );
  CFD2QXL \reg_mem_reg[5][9]  ( .D(n1206), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][9] ) );
  CFD2QXL \reg_mem_reg[5][10]  ( .D(n1205), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][10] ) );
  CFD2QXL \reg_mem_reg[5][11]  ( .D(n1204), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][11] ) );
  CFD2QXL \reg_mem_reg[5][12]  ( .D(n1203), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][12] ) );
  CFD2QXL \reg_mem_reg[4][11]  ( .D(n1236), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][11] ) );
  CFD2QXL \reg_mem_reg[4][12]  ( .D(n1235), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][12] ) );
  CFD2QXL \reg_mem_reg[3][0]  ( .D(n1279), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][0] ) );
  CFD2QXL \reg_mem_reg[3][2]  ( .D(n1277), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][2] ) );
  CFD2QXL \reg_mem_reg[3][3]  ( .D(n1276), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][3] ) );
  CFD2QXL \reg_mem_reg[3][4]  ( .D(n1275), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][4] ) );
  CFD2QXL \reg_mem_reg[3][5]  ( .D(n1274), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][5] ) );
  CFD2QXL \reg_mem_reg[3][6]  ( .D(n1273), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][6] ) );
  CFD2QXL \reg_mem_reg[3][7]  ( .D(n1272), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][7] ) );
  CFD2QXL \reg_mem_reg[3][8]  ( .D(n1271), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][8] ) );
  CFD2QXL \reg_mem_reg[3][9]  ( .D(n1270), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][9] ) );
  CFD2QXL \reg_mem_reg[3][10]  ( .D(n1269), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][10] ) );
  CFD2QXL \reg_mem_reg[31][0]  ( .D(n383), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][0] ) );
  CFD2QXL \reg_mem_reg[31][1]  ( .D(n382), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][1] ) );
  CFD2QXL \reg_mem_reg[31][2]  ( .D(n381), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][2] ) );
  CFD2QXL \reg_mem_reg[31][3]  ( .D(n380), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][3] ) );
  CFD2QXL \reg_mem_reg[31][4]  ( .D(n379), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][4] ) );
  CFD2QXL \reg_mem_reg[31][6]  ( .D(n377), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][6] ) );
  CFD2QXL \reg_mem_reg[31][8]  ( .D(n375), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][8] ) );
  CFD2QXL \reg_mem_reg[31][9]  ( .D(n374), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][9] ) );
  CFD2QXL \reg_mem_reg[31][10]  ( .D(n373), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][10] ) );
  CFD2QXL \reg_mem_reg[31][11]  ( .D(n372), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][11] ) );
  CFD2QXL \reg_mem_reg[31][12]  ( .D(n371), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][12] ) );
  CFD2QXL \reg_mem_reg[31][13]  ( .D(n370), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][13] ) );
  CFD2QXL \reg_mem_reg[31][14]  ( .D(n369), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][14] ) );
  CFD2QXL \reg_mem_reg[31][16]  ( .D(n367), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][16] ) );
  CFD2QXL \reg_mem_reg[31][17]  ( .D(n366), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][17] ) );
  CFD2QXL \reg_mem_reg[31][18]  ( .D(n365), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][18] ) );
  CFD2QXL \reg_mem_reg[31][19]  ( .D(n364), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][19] ) );
  CFD2QXL \reg_mem_reg[31][24]  ( .D(n359), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][24] ) );
  CFD2QXL \reg_mem_reg[31][27]  ( .D(n356), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][27] ) );
  CFD2QXL \reg_mem_reg[31][28]  ( .D(n355), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][28] ) );
  CFD2QXL \reg_mem_reg[31][30]  ( .D(n353), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][30] ) );
  CFD2QXL \reg_mem_reg[7][0]  ( .D(n1151), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][0] ) );
  CFD2QXL \reg_mem_reg[7][1]  ( .D(n1150), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][1] ) );
  CFD2QXL \reg_mem_reg[7][2]  ( .D(n1149), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][2] ) );
  CFD2QXL \reg_mem_reg[7][3]  ( .D(n1148), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][3] ) );
  CFD2QXL \reg_mem_reg[7][4]  ( .D(n1147), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][4] ) );
  CFD2QXL \reg_mem_reg[7][5]  ( .D(n1146), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][5] ) );
  CFD2QXL \reg_mem_reg[7][6]  ( .D(n1145), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][6] ) );
  CFD2QXL \reg_mem_reg[7][7]  ( .D(n1144), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][7] ) );
  CFD2QXL \reg_mem_reg[7][8]  ( .D(n1143), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][8] ) );
  CFD2QXL \reg_mem_reg[7][9]  ( .D(n1142), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][9] ) );
  CFD2QXL \reg_mem_reg[7][10]  ( .D(n1141), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][10] ) );
  CFD2QXL \reg_mem_reg[7][11]  ( .D(n1140), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][11] ) );
  CFD2QXL \reg_mem_reg[7][12]  ( .D(n1139), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][12] ) );
  CFD2QXL \reg_mem_reg[30][12]  ( .D(n403), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][12] ) );
  CFD2QXL \reg_mem_reg[30][13]  ( .D(n402), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][13] ) );
  CFD2QXL \reg_mem_reg[30][14]  ( .D(n401), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][14] ) );
  CFD2QXL \reg_mem_reg[30][16]  ( .D(n399), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][16] ) );
  CFD2QXL \reg_mem_reg[30][17]  ( .D(n398), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][17] ) );
  CFD2QXL \reg_mem_reg[30][18]  ( .D(n397), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][18] ) );
  CFD2QXL \reg_mem_reg[30][19]  ( .D(n396), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][19] ) );
  CFD2QXL \reg_mem_reg[30][24]  ( .D(n391), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][24] ) );
  CFD2QXL \reg_mem_reg[30][27]  ( .D(n388), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][27] ) );
  CFD2QXL \reg_mem_reg[30][28]  ( .D(n387), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][28] ) );
  CFD2QXL \reg_mem_reg[30][30]  ( .D(n385), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][30] ) );
  CFD2QXL \reg_mem_reg[6][1]  ( .D(n1182), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][1] ) );
  CFD2QXL \reg_mem_reg[6][11]  ( .D(n1172), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][11] ) );
  CFD2QXL \reg_mem_reg[6][12]  ( .D(n1171), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][12] ) );
  CFD2QXL \reg_mem_reg[9][0]  ( .D(n1087), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][0] ) );
  CFD2QXL \reg_mem_reg[9][2]  ( .D(n1085), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][2] ) );
  CFD2QXL \reg_mem_reg[9][3]  ( .D(n1084), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][3] ) );
  CFD2QXL \reg_mem_reg[9][4]  ( .D(n1083), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][4] ) );
  CFD2QXL \reg_mem_reg[9][5]  ( .D(n1082), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][5] ) );
  CFD2QXL \reg_mem_reg[9][6]  ( .D(n1081), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][6] ) );
  CFD2QXL \reg_mem_reg[9][7]  ( .D(n1080), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][7] ) );
  CFD2QXL \reg_mem_reg[9][8]  ( .D(n1079), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][8] ) );
  CFD2QXL \reg_mem_reg[9][9]  ( .D(n1078), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][9] ) );
  CFD2QXL \reg_mem_reg[9][10]  ( .D(n1077), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][10] ) );
  CFD2QXL \reg_mem_reg[9][13]  ( .D(n1074), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][13] ) );
  CFD2QXL \reg_mem_reg[9][14]  ( .D(n1073), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][14] ) );
  CFD2QXL \reg_mem_reg[9][16]  ( .D(n1071), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][16] ) );
  CFD2QXL \reg_mem_reg[9][17]  ( .D(n1070), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][17] ) );
  CFD2QXL \reg_mem_reg[9][19]  ( .D(n1068), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][19] ) );
  CFD2QXL \reg_mem_reg[1][0]  ( .D(n1343), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][0] ) );
  CFD2QXL \reg_mem_reg[1][2]  ( .D(n1341), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][2] ) );
  CFD2QXL \reg_mem_reg[1][3]  ( .D(n1340), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][3] ) );
  CFD2QXL \reg_mem_reg[1][4]  ( .D(n1339), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][4] ) );
  CFD2QXL \reg_mem_reg[1][5]  ( .D(n1338), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][5] ) );
  CFD2QXL \reg_mem_reg[1][6]  ( .D(n1337), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][6] ) );
  CFD2QXL \reg_mem_reg[1][7]  ( .D(n1336), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][7] ) );
  CFD2QXL \reg_mem_reg[1][9]  ( .D(n1334), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][9] ) );
  CFD2QXL \reg_mem_reg[1][10]  ( .D(n1333), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][10] ) );
  CFD2QXL \reg_mem_reg[8][13]  ( .D(n1106), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][13] ) );
  CFD2QXL \reg_mem_reg[8][14]  ( .D(n1105), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][14] ) );
  CFD2QXL \reg_mem_reg[8][16]  ( .D(n1103), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][16] ) );
  CFD2QXL \reg_mem_reg[8][17]  ( .D(n1102), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][17] ) );
  CFD2QXL \reg_mem_reg[8][19]  ( .D(n1100), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][19] ) );
  CFD2QXL \reg_mem_reg[5][13]  ( .D(n1202), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][13] ) );
  CFD2QXL \reg_mem_reg[5][14]  ( .D(n1201), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][14] ) );
  CFD2QXL \reg_mem_reg[5][16]  ( .D(n1199), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][16] ) );
  CFD2QXL \reg_mem_reg[5][17]  ( .D(n1198), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][17] ) );
  CFD2QXL \reg_mem_reg[5][18]  ( .D(n1197), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][18] ) );
  CFD2QXL \reg_mem_reg[5][19]  ( .D(n1196), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][19] ) );
  CFD2QXL \reg_mem_reg[5][24]  ( .D(n1191), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][24] ) );
  CFD2QXL \reg_mem_reg[5][27]  ( .D(n1188), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][27] ) );
  CFD2QXL \reg_mem_reg[5][28]  ( .D(n1187), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][28] ) );
  CFD2QXL \reg_mem_reg[5][30]  ( .D(n1185), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][30] ) );
  CFD2QXL \reg_mem_reg[5][31]  ( .D(n1184), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][31] ) );
  CFD2QXL \reg_mem_reg[4][3]  ( .D(n1244), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][3] ) );
  CFD2QXL \reg_mem_reg[4][4]  ( .D(n1243), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][4] ) );
  CFD2QXL \reg_mem_reg[4][5]  ( .D(n1242), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][5] ) );
  CFD2QXL \reg_mem_reg[4][6]  ( .D(n1241), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][6] ) );
  CFD2QXL \reg_mem_reg[4][7]  ( .D(n1240), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][7] ) );
  CFD2QXL \reg_mem_reg[4][9]  ( .D(n1238), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][9] ) );
  CFD2QXL \reg_mem_reg[4][10]  ( .D(n1237), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][10] ) );
  CFD2QXL \reg_mem_reg[4][13]  ( .D(n1234), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][13] ) );
  CFD2QXL \reg_mem_reg[4][14]  ( .D(n1233), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][14] ) );
  CFD2QXL \reg_mem_reg[4][15]  ( .D(n1232), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][15] ) );
  CFD2QXL \reg_mem_reg[4][16]  ( .D(n1231), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][16] ) );
  CFD2QXL \reg_mem_reg[4][17]  ( .D(n1230), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][17] ) );
  CFD2QXL \reg_mem_reg[4][18]  ( .D(n1229), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][18] ) );
  CFD2QXL \reg_mem_reg[4][19]  ( .D(n1228), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][19] ) );
  CFD2QXL \reg_mem_reg[4][21]  ( .D(n1226), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][21] ) );
  CFD2QXL \reg_mem_reg[4][24]  ( .D(n1223), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][24] ) );
  CFD2QXL \reg_mem_reg[4][27]  ( .D(n1220), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][27] ) );
  CFD2QXL \reg_mem_reg[4][28]  ( .D(n1219), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][28] ) );
  CFD2QXL \reg_mem_reg[4][30]  ( .D(n1217), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][30] ) );
  CFD2QXL \reg_mem_reg[3][1]  ( .D(n1278), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][1] ) );
  CFD2QXL \reg_mem_reg[3][11]  ( .D(n1268), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][11] ) );
  CFD2QXL \reg_mem_reg[3][12]  ( .D(n1267), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][12] ) );
  CFD2QXL \reg_mem_reg[3][13]  ( .D(n1266), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][13] ) );
  CFD2QXL \reg_mem_reg[3][14]  ( .D(n1265), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][14] ) );
  CFD2QXL \reg_mem_reg[3][16]  ( .D(n1263), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][16] ) );
  CFD2QXL \reg_mem_reg[3][17]  ( .D(n1262), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][17] ) );
  CFD2QXL \reg_mem_reg[3][18]  ( .D(n1261), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][18] ) );
  CFD2QXL \reg_mem_reg[3][19]  ( .D(n1260), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][19] ) );
  CFD2QXL \reg_mem_reg[3][24]  ( .D(n1255), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][24] ) );
  CFD2QXL \reg_mem_reg[3][27]  ( .D(n1252), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][27] ) );
  CFD2QXL \reg_mem_reg[3][28]  ( .D(n1251), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][28] ) );
  CFD2QXL \reg_mem_reg[3][30]  ( .D(n1249), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][30] ) );
  CFD2QXL \reg_mem_reg[2][0]  ( .D(n1311), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][0] ) );
  CFD2QXL \reg_mem_reg[2][1]  ( .D(n1310), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][1] ) );
  CFD2QXL \reg_mem_reg[2][2]  ( .D(n1309), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][2] ) );
  CFD2QXL \reg_mem_reg[2][3]  ( .D(n1308), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][3] ) );
  CFD2QXL \reg_mem_reg[2][4]  ( .D(n1307), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][4] ) );
  CFD2QXL \reg_mem_reg[2][5]  ( .D(n1306), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][5] ) );
  CFD2QXL \reg_mem_reg[2][6]  ( .D(n1305), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][6] ) );
  CFD2QXL \reg_mem_reg[2][7]  ( .D(n1304), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][7] ) );
  CFD2QXL \reg_mem_reg[2][8]  ( .D(n1303), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][8] ) );
  CFD2QXL \reg_mem_reg[2][9]  ( .D(n1302), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][9] ) );
  CFD2QXL \reg_mem_reg[2][10]  ( .D(n1301), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][10] ) );
  CFD2QXL \reg_mem_reg[2][11]  ( .D(n1300), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][11] ) );
  CFD2QXL \reg_mem_reg[2][12]  ( .D(n1299), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][12] ) );
  CFD2QXL \reg_mem_reg[2][13]  ( .D(n1298), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][13] ) );
  CFD2QXL \reg_mem_reg[2][14]  ( .D(n1297), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][14] ) );
  CFD2QXL \reg_mem_reg[2][16]  ( .D(n1295), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][16] ) );
  CFD2QXL \reg_mem_reg[2][17]  ( .D(n1294), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][17] ) );
  CFD2QXL \reg_mem_reg[2][18]  ( .D(n1293), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][18] ) );
  CFD2QXL \reg_mem_reg[2][19]  ( .D(n1292), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][19] ) );
  CFD2QXL \reg_mem_reg[2][24]  ( .D(n1287), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][24] ) );
  CFD2QXL \reg_mem_reg[2][27]  ( .D(n1284), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][27] ) );
  CFD2QXL \reg_mem_reg[2][28]  ( .D(n1283), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][28] ) );
  CFD2QXL \reg_mem_reg[2][30]  ( .D(n1281), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][30] ) );
  CFD2QXL \reg_mem_reg[7][13]  ( .D(n1138), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][13] ) );
  CFD2QXL \reg_mem_reg[7][14]  ( .D(n1137), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][14] ) );
  CFD2QXL \reg_mem_reg[7][16]  ( .D(n1135), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][16] ) );
  CFD2QXL \reg_mem_reg[7][17]  ( .D(n1134), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][17] ) );
  CFD2QXL \reg_mem_reg[7][18]  ( .D(n1133), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][18] ) );
  CFD2QXL \reg_mem_reg[7][19]  ( .D(n1132), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][19] ) );
  CFD2QXL \reg_mem_reg[7][24]  ( .D(n1127), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][24] ) );
  CFD2QXL \reg_mem_reg[7][27]  ( .D(n1124), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][27] ) );
  CFD2QXL \reg_mem_reg[7][28]  ( .D(n1123), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][28] ) );
  CFD2QXL \reg_mem_reg[7][30]  ( .D(n1121), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][30] ) );
  CFD2QXL \reg_mem_reg[7][31]  ( .D(n1120), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][31] ) );
  CFD2QXL \reg_mem_reg[30][0]  ( .D(n415), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][0] ) );
  CFD2QXL \reg_mem_reg[30][1]  ( .D(n414), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][1] ) );
  CFD2QXL \reg_mem_reg[30][2]  ( .D(n413), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][2] ) );
  CFD2QXL \reg_mem_reg[30][3]  ( .D(n412), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][3] ) );
  CFD2QXL \reg_mem_reg[30][4]  ( .D(n411), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][4] ) );
  CFD2QXL \reg_mem_reg[30][5]  ( .D(n410), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][5] ) );
  CFD2QXL \reg_mem_reg[30][6]  ( .D(n409), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][6] ) );
  CFD2QXL \reg_mem_reg[30][7]  ( .D(n408), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][7] ) );
  CFD2QXL \reg_mem_reg[30][8]  ( .D(n407), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][8] ) );
  CFD2QXL \reg_mem_reg[30][9]  ( .D(n406), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][9] ) );
  CFD2QXL \reg_mem_reg[30][10]  ( .D(n405), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][10] ) );
  CFD2QXL \reg_mem_reg[30][11]  ( .D(n404), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][11] ) );
  CFD2QXL \reg_mem_reg[6][0]  ( .D(n1183), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][0] ) );
  CFD2QXL \reg_mem_reg[6][2]  ( .D(n1181), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][2] ) );
  CFD2QXL \reg_mem_reg[6][3]  ( .D(n1180), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][3] ) );
  CFD2QXL \reg_mem_reg[6][4]  ( .D(n1179), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][4] ) );
  CFD2QXL \reg_mem_reg[6][5]  ( .D(n1178), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][5] ) );
  CFD2QXL \reg_mem_reg[6][6]  ( .D(n1177), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][6] ) );
  CFD2QXL \reg_mem_reg[6][7]  ( .D(n1176), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][7] ) );
  CFD2QXL \reg_mem_reg[6][8]  ( .D(n1175), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][8] ) );
  CFD2QXL \reg_mem_reg[6][9]  ( .D(n1174), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][9] ) );
  CFD2QXL \reg_mem_reg[6][10]  ( .D(n1173), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][10] ) );
  CFD2QXL \reg_mem_reg[6][13]  ( .D(n1170), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][13] ) );
  CFD2QXL \reg_mem_reg[6][14]  ( .D(n1169), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][14] ) );
  CFD2QXL \reg_mem_reg[6][15]  ( .D(n1168), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][15] ) );
  CFD2QXL \reg_mem_reg[6][16]  ( .D(n1167), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][16] ) );
  CFD2QXL \reg_mem_reg[6][17]  ( .D(n1166), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][17] ) );
  CFD2QXL \reg_mem_reg[6][18]  ( .D(n1165), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][18] ) );
  CFD2QXL \reg_mem_reg[6][19]  ( .D(n1164), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][19] ) );
  CFD2QXL \reg_mem_reg[6][21]  ( .D(n1162), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][21] ) );
  CFD2QXL \reg_mem_reg[6][24]  ( .D(n1159), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][24] ) );
  CFD2QXL \reg_mem_reg[6][27]  ( .D(n1156), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][27] ) );
  CFD2QXL \reg_mem_reg[6][28]  ( .D(n1155), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][28] ) );
  CFD2QXL \reg_mem_reg[6][30]  ( .D(n1153), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][30] ) );
  CFD2QXL \reg_mem_reg[9][1]  ( .D(n1086), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][1] ) );
  CFD2QXL \reg_mem_reg[9][11]  ( .D(n1076), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][11] ) );
  CFD2QXL \reg_mem_reg[9][12]  ( .D(n1075), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][12] ) );
  CFD2QXL \reg_mem_reg[9][18]  ( .D(n1069), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][18] ) );
  CFD2QXL \reg_mem_reg[9][24]  ( .D(n1063), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][24] ) );
  CFD2QXL \reg_mem_reg[9][27]  ( .D(n1060), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][27] ) );
  CFD2QXL \reg_mem_reg[9][28]  ( .D(n1059), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][28] ) );
  CFD2QXL \reg_mem_reg[9][30]  ( .D(n1057), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][30] ) );
  CFD2QXL \reg_mem_reg[9][31]  ( .D(n1056), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][31] ) );
  CFD2QXL \reg_mem_reg[1][1]  ( .D(n1342), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][1] ) );
  CFD2QXL \reg_mem_reg[1][11]  ( .D(n1332), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][11] ) );
  CFD2QXL \reg_mem_reg[1][12]  ( .D(n1331), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][12] ) );
  CFD2QXL \reg_mem_reg[1][13]  ( .D(n1330), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][13] ) );
  CFD2QXL \reg_mem_reg[1][14]  ( .D(n1329), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][14] ) );
  CFD2QXL \reg_mem_reg[1][16]  ( .D(n1327), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][16] ) );
  CFD2QXL \reg_mem_reg[1][17]  ( .D(n1326), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][17] ) );
  CFD2QXL \reg_mem_reg[1][18]  ( .D(n1325), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][18] ) );
  CFD2QXL \reg_mem_reg[1][19]  ( .D(n1324), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][19] ) );
  CFD2QXL \reg_mem_reg[1][24]  ( .D(n1319), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][24] ) );
  CFD2QXL \reg_mem_reg[1][27]  ( .D(n1316), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][27] ) );
  CFD2QXL \reg_mem_reg[1][28]  ( .D(n1315), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][28] ) );
  CFD2QXL \reg_mem_reg[1][30]  ( .D(n1313), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][30] ) );
  CFD2QXL \reg_mem_reg[8][0]  ( .D(n1119), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][0] ) );
  CFD2QXL \reg_mem_reg[8][1]  ( .D(n1118), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][1] ) );
  CFD2QXL \reg_mem_reg[8][2]  ( .D(n1117), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][2] ) );
  CFD2QXL \reg_mem_reg[8][3]  ( .D(n1116), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][3] ) );
  CFD2QXL \reg_mem_reg[8][4]  ( .D(n1115), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][4] ) );
  CFD2QXL \reg_mem_reg[8][5]  ( .D(n1114), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][5] ) );
  CFD2QXL \reg_mem_reg[8][6]  ( .D(n1113), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][6] ) );
  CFD2QXL \reg_mem_reg[8][7]  ( .D(n1112), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][7] ) );
  CFD2QXL \reg_mem_reg[8][8]  ( .D(n1111), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][8] ) );
  CFD2QXL \reg_mem_reg[8][9]  ( .D(n1110), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][9] ) );
  CFD2QXL \reg_mem_reg[8][10]  ( .D(n1109), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][10] ) );
  CFD2QXL \reg_mem_reg[8][11]  ( .D(n1108), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][11] ) );
  CFD2QXL \reg_mem_reg[8][12]  ( .D(n1107), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][12] ) );
  CFD2QXL \reg_mem_reg[8][18]  ( .D(n1101), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][18] ) );
  CFD2QXL \reg_mem_reg[8][24]  ( .D(n1095), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][24] ) );
  CFD2QXL \reg_mem_reg[8][27]  ( .D(n1092), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][27] ) );
  CFD2QXL \reg_mem_reg[8][28]  ( .D(n1091), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][28] ) );
  CFD2QXL \reg_mem_reg[8][30]  ( .D(n1089), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][30] ) );
  CFD2QXL \reg_mem_reg[0][0]  ( .D(n1375), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][0] ) );
  CFD2QXL \reg_mem_reg[0][1]  ( .D(n1374), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][1] ) );
  CFD2QXL \reg_mem_reg[0][2]  ( .D(n1373), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][2] ) );
  CFD2QXL \reg_mem_reg[0][3]  ( .D(n1372), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][3] ) );
  CFD2QXL \reg_mem_reg[0][4]  ( .D(n1371), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][4] ) );
  CFD2QXL \reg_mem_reg[0][5]  ( .D(n1370), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][5] ) );
  CFD2QXL \reg_mem_reg[0][6]  ( .D(n1369), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][6] ) );
  CFD2QXL \reg_mem_reg[0][7]  ( .D(n1368), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][7] ) );
  CFD2QXL \reg_mem_reg[0][9]  ( .D(n1366), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][9] ) );
  CFD2QXL \reg_mem_reg[0][10]  ( .D(n1365), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][10] ) );
  CFD2QXL \reg_mem_reg[0][11]  ( .D(n1364), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][11] ) );
  CFD2QXL \reg_mem_reg[0][12]  ( .D(n1363), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][12] ) );
  CFD2QXL \reg_mem_reg[0][13]  ( .D(n1362), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][13] ) );
  CFD2QXL \reg_mem_reg[0][14]  ( .D(n1361), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][14] ) );
  CFD2QXL \reg_mem_reg[0][16]  ( .D(n1359), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][16] ) );
  CFD2QXL \reg_mem_reg[0][17]  ( .D(n1358), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][17] ) );
  CFD2QXL \reg_mem_reg[0][18]  ( .D(n1357), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][18] ) );
  CFD2QXL \reg_mem_reg[0][19]  ( .D(n1356), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][19] ) );
  CFD2QXL \reg_mem_reg[0][24]  ( .D(n1351), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][24] ) );
  CFD2QXL \reg_mem_reg[0][27]  ( .D(n1348), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][27] ) );
  CFD2QXL \reg_mem_reg[0][28]  ( .D(n1347), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][28] ) );
  CFD2QXL \reg_mem_reg[0][30]  ( .D(n1345), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][30] ) );
  CFD2QXL \opcode_mem_reg[0]  ( .D(n1843), .CP(clk), .CD(rst), .Q(
        opcode_mem[0]) );
  CFD2QXL \opcode_mem_reg[1]  ( .D(n1844), .CP(clk), .CD(rst), .Q(
        opcode_mem[1]) );
  CFD2QXL \prog_count_reg[6]  ( .D(prog_count_c[6]), .CP(clk), .CD(rst), .Q(
        prog_count_o[6]) );
  CFD2QXL \prog_count_reg[5]  ( .D(prog_count_c[5]), .CP(clk), .CD(rst), .Q(
        prog_count_o[5]) );
  CFD1QXL \reg_mem_reg[21][22]  ( .D(n681), .CP(clk), .Q(\reg_mem[21][22] ) );
  CFD1QXL \reg_mem_reg[21][25]  ( .D(n678), .CP(clk), .Q(\reg_mem[21][25] ) );
  CFD1QXL \reg_mem_reg[21][26]  ( .D(n677), .CP(clk), .Q(\reg_mem[21][26] ) );
  CFD1QXL \reg_mem_reg[13][22]  ( .D(n937), .CP(clk), .Q(\reg_mem[13][22] ) );
  CFD1QXL \reg_mem_reg[13][25]  ( .D(n934), .CP(clk), .Q(\reg_mem[13][25] ) );
  CFD1QXL \reg_mem_reg[13][26]  ( .D(n933), .CP(clk), .Q(\reg_mem[13][26] ) );
  CFD1QXL \reg_mem_reg[28][22]  ( .D(n457), .CP(clk), .Q(\reg_mem[28][22] ) );
  CFD1QXL \reg_mem_reg[28][25]  ( .D(n454), .CP(clk), .Q(\reg_mem[28][25] ) );
  CFD1QXL \reg_mem_reg[28][26]  ( .D(n453), .CP(clk), .Q(\reg_mem[28][26] ) );
  CFD1QXL \reg_mem_reg[20][22]  ( .D(n713), .CP(clk), .Q(\reg_mem[20][22] ) );
  CFD1QXL \reg_mem_reg[20][25]  ( .D(n710), .CP(clk), .Q(\reg_mem[20][25] ) );
  CFD1QXL \reg_mem_reg[20][26]  ( .D(n709), .CP(clk), .Q(\reg_mem[20][26] ) );
  CFD1QXL \reg_mem_reg[12][22]  ( .D(n969), .CP(clk), .Q(\reg_mem[12][22] ) );
  CFD1QXL \reg_mem_reg[12][25]  ( .D(n966), .CP(clk), .Q(\reg_mem[12][25] ) );
  CFD1QXL \reg_mem_reg[12][26]  ( .D(n965), .CP(clk), .Q(\reg_mem[12][26] ) );
  CFD1QXL \reg_mem_reg[27][22]  ( .D(n489), .CP(clk), .Q(\reg_mem[27][22] ) );
  CFD1QXL \reg_mem_reg[27][25]  ( .D(n486), .CP(clk), .Q(\reg_mem[27][25] ) );
  CFD1QXL \reg_mem_reg[27][26]  ( .D(n485), .CP(clk), .Q(\reg_mem[27][26] ) );
  CFD1QXL \reg_mem_reg[19][22]  ( .D(n745), .CP(clk), .Q(\reg_mem[19][22] ) );
  CFD1QXL \reg_mem_reg[19][25]  ( .D(n742), .CP(clk), .Q(\reg_mem[19][25] ) );
  CFD1QXL \reg_mem_reg[19][26]  ( .D(n741), .CP(clk), .Q(\reg_mem[19][26] ) );
  CFD1QXL \reg_mem_reg[11][22]  ( .D(n1001), .CP(clk), .Q(\reg_mem[11][22] )
         );
  CFD1QXL \reg_mem_reg[11][25]  ( .D(n998), .CP(clk), .Q(\reg_mem[11][25] ) );
  CFD1QXL \reg_mem_reg[11][26]  ( .D(n997), .CP(clk), .Q(\reg_mem[11][26] ) );
  CFD1QXL \reg_mem_reg[26][22]  ( .D(n521), .CP(clk), .Q(\reg_mem[26][22] ) );
  CFD1QXL \reg_mem_reg[26][25]  ( .D(n518), .CP(clk), .Q(\reg_mem[26][25] ) );
  CFD1QXL \reg_mem_reg[18][22]  ( .D(n777), .CP(clk), .Q(\reg_mem[18][22] ) );
  CFD1QXL \reg_mem_reg[18][25]  ( .D(n774), .CP(clk), .Q(\reg_mem[18][25] ) );
  CFD1QXL \reg_mem_reg[18][26]  ( .D(n773), .CP(clk), .Q(\reg_mem[18][26] ) );
  CFD1QXL \reg_mem_reg[18][31]  ( .D(n768), .CP(clk), .Q(\reg_mem[18][31] ) );
  CFD1QXL \reg_mem_reg[10][22]  ( .D(n1033), .CP(clk), .Q(\reg_mem[10][22] )
         );
  CFD1QXL \reg_mem_reg[10][25]  ( .D(n1030), .CP(clk), .Q(\reg_mem[10][25] )
         );
  CFD1QXL \reg_mem_reg[23][22]  ( .D(n617), .CP(clk), .Q(\reg_mem[23][22] ) );
  CFD1QXL \reg_mem_reg[23][25]  ( .D(n614), .CP(clk), .Q(\reg_mem[23][25] ) );
  CFD1QXL \reg_mem_reg[23][26]  ( .D(n613), .CP(clk), .Q(\reg_mem[23][26] ) );
  CFD1QXL \reg_mem_reg[15][22]  ( .D(n873), .CP(clk), .Q(\reg_mem[15][22] ) );
  CFD1QXL \reg_mem_reg[15][25]  ( .D(n870), .CP(clk), .Q(\reg_mem[15][25] ) );
  CFD1QXL \reg_mem_reg[15][26]  ( .D(n869), .CP(clk), .Q(\reg_mem[15][26] ) );
  CFD1QXL \reg_mem_reg[22][22]  ( .D(n649), .CP(clk), .Q(\reg_mem[22][22] ) );
  CFD1QXL \reg_mem_reg[22][25]  ( .D(n646), .CP(clk), .Q(\reg_mem[22][25] ) );
  CFD1QXL \reg_mem_reg[22][26]  ( .D(n645), .CP(clk), .Q(\reg_mem[22][26] ) );
  CFD1QXL \reg_mem_reg[14][22]  ( .D(n905), .CP(clk), .Q(\reg_mem[14][22] ) );
  CFD1QXL \reg_mem_reg[14][25]  ( .D(n902), .CP(clk), .Q(\reg_mem[14][25] ) );
  CFD1QXL \reg_mem_reg[14][26]  ( .D(n901), .CP(clk), .Q(\reg_mem[14][26] ) );
  CFD1QXL \reg_mem_reg[25][22]  ( .D(n553), .CP(clk), .Q(\reg_mem[25][22] ) );
  CFD1QXL \reg_mem_reg[25][25]  ( .D(n550), .CP(clk), .Q(\reg_mem[25][25] ) );
  CFD1QXL \reg_mem_reg[25][26]  ( .D(n549), .CP(clk), .Q(\reg_mem[25][26] ) );
  CFD1QXL \reg_mem_reg[17][22]  ( .D(n809), .CP(clk), .Q(\reg_mem[17][22] ) );
  CFD1QXL \reg_mem_reg[17][25]  ( .D(n806), .CP(clk), .Q(\reg_mem[17][25] ) );
  CFD1QXL \reg_mem_reg[17][26]  ( .D(n805), .CP(clk), .Q(\reg_mem[17][26] ) );
  CFD1QXL \reg_mem_reg[24][22]  ( .D(n585), .CP(clk), .Q(\reg_mem[24][22] ) );
  CFD1QXL \reg_mem_reg[24][26]  ( .D(n581), .CP(clk), .Q(\reg_mem[24][26] ) );
  CFD1QXL \reg_mem_reg[16][22]  ( .D(n841), .CP(clk), .Q(\reg_mem[16][22] ) );
  CFD1QXL \reg_mem_reg[16][25]  ( .D(n838), .CP(clk), .Q(\reg_mem[16][25] ) );
  CFD1QXL \reg_mem_reg[16][26]  ( .D(n837), .CP(clk), .Q(\reg_mem[16][26] ) );
  CFD1QXL \reg_mem_reg[16][31]  ( .D(n832), .CP(clk), .Q(\reg_mem[16][31] ) );
  CFD1QXL \reg_mem_reg[13][20]  ( .D(n939), .CP(clk), .Q(\reg_mem[13][20] ) );
  CFD1QXL \reg_mem_reg[13][23]  ( .D(n936), .CP(clk), .Q(\reg_mem[13][23] ) );
  CFD1QXL \reg_mem_reg[28][20]  ( .D(n459), .CP(clk), .Q(\reg_mem[28][20] ) );
  CFD1QXL \reg_mem_reg[28][23]  ( .D(n456), .CP(clk), .Q(\reg_mem[28][23] ) );
  CFD1QXL \reg_mem_reg[12][20]  ( .D(n971), .CP(clk), .Q(\reg_mem[12][20] ) );
  CFD1QXL \reg_mem_reg[12][23]  ( .D(n968), .CP(clk), .Q(\reg_mem[12][23] ) );
  CFD1QXL \reg_mem_reg[27][20]  ( .D(n491), .CP(clk), .Q(\reg_mem[27][20] ) );
  CFD1QXL \reg_mem_reg[27][23]  ( .D(n488), .CP(clk), .Q(\reg_mem[27][23] ) );
  CFD1QXL \reg_mem_reg[11][20]  ( .D(n1003), .CP(clk), .Q(\reg_mem[11][20] )
         );
  CFD1QXL \reg_mem_reg[11][23]  ( .D(n1000), .CP(clk), .Q(\reg_mem[11][23] )
         );
  CFD1QXL \reg_mem_reg[26][20]  ( .D(n523), .CP(clk), .Q(\reg_mem[26][20] ) );
  CFD1QXL \reg_mem_reg[26][23]  ( .D(n520), .CP(clk), .Q(\reg_mem[26][23] ) );
  CFD1QXL \reg_mem_reg[10][20]  ( .D(n1035), .CP(clk), .Q(\reg_mem[10][20] )
         );
  CFD1QXL \reg_mem_reg[10][23]  ( .D(n1032), .CP(clk), .Q(\reg_mem[10][23] )
         );
  CFD1QXL \reg_mem_reg[15][20]  ( .D(n875), .CP(clk), .Q(\reg_mem[15][20] ) );
  CFD1QXL \reg_mem_reg[15][23]  ( .D(n872), .CP(clk), .Q(\reg_mem[15][23] ) );
  CFD1QXL \reg_mem_reg[14][20]  ( .D(n907), .CP(clk), .Q(\reg_mem[14][20] ) );
  CFD1QXL \reg_mem_reg[14][23]  ( .D(n904), .CP(clk), .Q(\reg_mem[14][23] ) );
  CFD1QXL \reg_mem_reg[25][20]  ( .D(n555), .CP(clk), .Q(\reg_mem[25][20] ) );
  CFD1QXL \reg_mem_reg[25][23]  ( .D(n552), .CP(clk), .Q(\reg_mem[25][23] ) );
  CFD1QXL \reg_mem_reg[17][29]  ( .D(n802), .CP(clk), .Q(\reg_mem[17][29] ) );
  CFD1QXL \reg_mem_reg[24][20]  ( .D(n587), .CP(clk), .Q(\reg_mem[24][20] ) );
  CFD1QXL \reg_mem_reg[24][23]  ( .D(n584), .CP(clk), .Q(\reg_mem[24][23] ) );
  CFD1QXL \reg_mem_reg[21][20]  ( .D(n683), .CP(clk), .Q(\reg_mem[21][20] ) );
  CFD1QXL \reg_mem_reg[21][23]  ( .D(n680), .CP(clk), .Q(\reg_mem[21][23] ) );
  CFD1QXL \reg_mem_reg[20][20]  ( .D(n715), .CP(clk), .Q(\reg_mem[20][20] ) );
  CFD1QXL \reg_mem_reg[20][23]  ( .D(n712), .CP(clk), .Q(\reg_mem[20][23] ) );
  CFD1QXL \reg_mem_reg[19][20]  ( .D(n747), .CP(clk), .Q(\reg_mem[19][20] ) );
  CFD1QXL \reg_mem_reg[19][23]  ( .D(n744), .CP(clk), .Q(\reg_mem[19][23] ) );
  CFD1QXL \reg_mem_reg[18][20]  ( .D(n779), .CP(clk), .Q(\reg_mem[18][20] ) );
  CFD1QXL \reg_mem_reg[18][23]  ( .D(n776), .CP(clk), .Q(\reg_mem[18][23] ) );
  CFD1QXL \reg_mem_reg[23][20]  ( .D(n619), .CP(clk), .Q(\reg_mem[23][20] ) );
  CFD1QXL \reg_mem_reg[22][20]  ( .D(n651), .CP(clk), .Q(\reg_mem[22][20] ) );
  CFD1QXL \reg_mem_reg[22][23]  ( .D(n648), .CP(clk), .Q(\reg_mem[22][23] ) );
  CFD1QXL \reg_mem_reg[17][20]  ( .D(n811), .CP(clk), .Q(\reg_mem[17][20] ) );
  CFD1QXL \reg_mem_reg[17][23]  ( .D(n808), .CP(clk), .Q(\reg_mem[17][23] ) );
  CFD1QXL \reg_mem_reg[16][20]  ( .D(n843), .CP(clk), .Q(\reg_mem[16][20] ) );
  CFD1QXL \reg_mem_reg[16][23]  ( .D(n840), .CP(clk), .Q(\reg_mem[16][23] ) );
  CFD2QX1 r_type_wb_reg ( .D(n1845), .CP(clk), .CD(rst), .Q(r_type_wb) );
  CFD2QXL \opcode_ext_ex_reg[10]  ( .D(opcode_ext_c[10]), .CP(clk), .CD(rst), 
        .Q(opcode_ext_ex[10]) );
  CFD2QXL \opcode_ext_ex_reg[7]  ( .D(opcode_ext_c[7]), .CP(clk), .CD(rst), 
        .Q(opcode_ext_ex[7]) );
  CFD2QXL \opcode_ext_ex_reg[1]  ( .D(opcode_ext_c[1]), .CP(clk), .CD(rst), 
        .Q(opcode_ext_ex[1]) );
  CFD1QXL \reg_mem_reg[18][29]  ( .D(n770), .CP(clk), .Q(\reg_mem[18][29] ) );
  CFD2QXL \opcode_ext_ex_reg[4]  ( .D(opcode_ext_c[4]), .CP(clk), .CD(rst), 
        .Q(opcode_ext_ex[4]) );
  CFD2QXL \opcode_ext_ex_reg[2]  ( .D(opcode_ext_c[2]), .CP(clk), .CD(rst), 
        .Q(opcode_ext_ex[2]) );
  CFD2QXL \regc_addr_wb_reg[4]  ( .D(n1848), .CP(clk), .CD(rst), .Q(
        regc_addr_wb[4]) );
  CFD2QXL \regc_addr_wb_reg[3]  ( .D(n1851), .CP(clk), .CD(rst), .Q(
        regc_addr_wb[3]) );
  CFD2QXL \regc_addr_wb_reg[1]  ( .D(n1854), .CP(clk), .CD(rst), .Q(
        regc_addr_wb[1]) );
  CFD2QXL \regc_addr_wb_reg[0]  ( .D(n1857), .CP(clk), .CD(rst), .Q(
        regc_addr_wb[0]) );
  CFD2QXL \regc_addr_wb_reg[2]  ( .D(n1860), .CP(clk), .CD(rst), .Q(
        regc_addr_wb[2]) );
  CFD2QXL \opcode_ext_ex_reg[8]  ( .D(opcode_ext_c[8]), .CP(clk), .CD(rst), 
        .Q(opcode_ext_ex[8]) );
  CFD2QXL \opcode_ext_ex_reg[5]  ( .D(opcode_ext_c[5]), .CP(clk), .CD(rst), 
        .Q(opcode_ext_ex[5]) );
  CFD2QXL \opcode_ext_ex_reg[9]  ( .D(opcode_ext_c[9]), .CP(clk), .CD(rst), 
        .Q(opcode_ext_ex[9]) );
  CFD2QXL \opcode_ext_ex_reg[6]  ( .D(opcode_ext_c[6]), .CP(clk), .CD(rst), 
        .Q(opcode_ext_ex[6]) );
  CFD2QXL \opcode_ext_ex_reg[3]  ( .D(opcode_ext_c[3]), .CP(clk), .CD(rst), 
        .Q(opcode_ext_ex[3]) );
  CFD2QXL \opcode_ext_ex_reg[0]  ( .D(opcode_ext_c[0]), .CP(clk), .CD(rst), 
        .Q(opcode_ext_ex[0]) );
  CFD2QXL \regb_addr_wb_reg[4]  ( .D(n1863), .CP(clk), .CD(rst), .Q(
        regb_addr_wb[4]) );
  CFD2QXL \regb_addr_wb_reg[3]  ( .D(n1866), .CP(clk), .CD(rst), .Q(
        regb_addr_wb[3]) );
  CFD2QXL \regb_addr_wb_reg[0]  ( .D(n1869), .CP(clk), .CD(rst), .Q(
        regb_addr_wb[0]) );
  CFD2QXL \regb_addr_wb_reg[2]  ( .D(n1872), .CP(clk), .CD(rst), .Q(
        regb_addr_wb[2]) );
  CFD2QXL \regb_addr_wb_reg[1]  ( .D(n1875), .CP(clk), .CD(rst), .Q(
        regb_addr_wb[1]) );
  CFD2QXL \regb_addr_reg[0]  ( .D(net87798), .CP(clk), .CD(rst), .Q(
        regb_addr[0]) );
  CFD2QXL \reg_mem_reg[29][21]  ( .D(n426), .CP(clk), .CD(rst), .Q(
        \reg_mem[29][21] ) );
  CFD2QXL \reg_mem_reg[29][22]  ( .D(n425), .CP(clk), .CD(rst), .Q(
        \reg_mem[29][22] ) );
  CFD2QXL \reg_mem_reg[29][25]  ( .D(n422), .CP(clk), .CD(rst), .Q(
        \reg_mem[29][25] ) );
  CFD2QXL \reg_mem_reg[29][26]  ( .D(n421), .CP(clk), .CD(rst), .Q(
        \reg_mem[29][26] ) );
  CFD2QXL \reg_mem_reg[5][22]  ( .D(n1193), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][22] ) );
  CFD2QXL \reg_mem_reg[5][25]  ( .D(n1190), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][25] ) );
  CFD2QXL \reg_mem_reg[5][26]  ( .D(n1189), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][26] ) );
  CFD2QXL \reg_mem_reg[4][22]  ( .D(n1225), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][22] ) );
  CFD2QXL \reg_mem_reg[4][25]  ( .D(n1222), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][25] ) );
  CFD2QXL \reg_mem_reg[4][26]  ( .D(n1221), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][26] ) );
  CFD2QXL \reg_mem_reg[4][31]  ( .D(n1216), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][31] ) );
  CFD2QXL \reg_mem_reg[3][15]  ( .D(n1264), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][15] ) );
  CFD2QXL \reg_mem_reg[3][21]  ( .D(n1258), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][21] ) );
  CFD2QXL \reg_mem_reg[3][22]  ( .D(n1257), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][22] ) );
  CFD2QXL \reg_mem_reg[3][25]  ( .D(n1254), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][25] ) );
  CFD2QXL \reg_mem_reg[3][26]  ( .D(n1253), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][26] ) );
  CFD2QXL \reg_mem_reg[2][22]  ( .D(n1289), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][22] ) );
  CFD2QXL \reg_mem_reg[2][25]  ( .D(n1286), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][25] ) );
  CFD2QXL \reg_mem_reg[2][26]  ( .D(n1285), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][26] ) );
  CFD2QXL \reg_mem_reg[2][31]  ( .D(n1280), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][31] ) );
  CFD2QXL \reg_mem_reg[31][22]  ( .D(n361), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][22] ) );
  CFD2QXL \reg_mem_reg[31][25]  ( .D(n358), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][25] ) );
  CFD2QXL \reg_mem_reg[31][26]  ( .D(n357), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][26] ) );
  CFD2QXL \reg_mem_reg[7][22]  ( .D(n1129), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][22] ) );
  CFD2QXL \reg_mem_reg[7][25]  ( .D(n1126), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][25] ) );
  CFD2QXL \reg_mem_reg[7][26]  ( .D(n1125), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][26] ) );
  CFD2QXL \reg_mem_reg[30][15]  ( .D(n400), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][15] ) );
  CFD2QXL \reg_mem_reg[30][21]  ( .D(n394), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][21] ) );
  CFD2QXL \reg_mem_reg[30][22]  ( .D(n393), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][22] ) );
  CFD2QXL \reg_mem_reg[30][25]  ( .D(n390), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][25] ) );
  CFD2QXL \reg_mem_reg[30][26]  ( .D(n389), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][26] ) );
  CFD2QXL \reg_mem_reg[6][22]  ( .D(n1161), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][22] ) );
  CFD2QXL \reg_mem_reg[6][25]  ( .D(n1158), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][25] ) );
  CFD2QXL \reg_mem_reg[6][26]  ( .D(n1157), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][26] ) );
  CFD2QXL \reg_mem_reg[6][31]  ( .D(n1152), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][31] ) );
  CFD2QXL \reg_mem_reg[9][22]  ( .D(n1065), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][22] ) );
  CFD2QXL \reg_mem_reg[9][25]  ( .D(n1062), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][25] ) );
  CFD2QXL \reg_mem_reg[9][26]  ( .D(n1061), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][26] ) );
  CFD2QXL \reg_mem_reg[1][15]  ( .D(n1328), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][15] ) );
  CFD2QXL \reg_mem_reg[1][21]  ( .D(n1322), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][21] ) );
  CFD2QXL \reg_mem_reg[1][22]  ( .D(n1321), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][22] ) );
  CFD2QXL \reg_mem_reg[1][25]  ( .D(n1318), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][25] ) );
  CFD2QXL \reg_mem_reg[1][26]  ( .D(n1317), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][26] ) );
  CFD2QXL \reg_mem_reg[8][15]  ( .D(n1104), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][15] ) );
  CFD2QXL \reg_mem_reg[8][21]  ( .D(n1098), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][21] ) );
  CFD2QXL \reg_mem_reg[8][22]  ( .D(n1097), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][22] ) );
  CFD2QXL \reg_mem_reg[8][26]  ( .D(n1093), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][26] ) );
  CFD2QXL \reg_mem_reg[0][22]  ( .D(n1353), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][22] ) );
  CFD2QXL \reg_mem_reg[0][25]  ( .D(n1350), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][25] ) );
  CFD2QXL \reg_mem_reg[0][26]  ( .D(n1349), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][26] ) );
  CFD2QXL \reg_mem_reg[0][31]  ( .D(n1344), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][31] ) );
  CFD2QXL \reg_mem_reg[4][8]  ( .D(n1877), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][8] ) );
  CFD2QXL \reg_mem_reg[5][8]  ( .D(n1207), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][8] ) );
  CFD2QXL \reg_mem_reg[29][20]  ( .D(n427), .CP(clk), .CD(rst), .Q(
        \reg_mem[29][20] ) );
  CFD2QXL \reg_mem_reg[29][23]  ( .D(n424), .CP(clk), .CD(rst), .Q(
        \reg_mem[29][23] ) );
  CFD2QXL \reg_mem_reg[29][29]  ( .D(n418), .CP(clk), .CD(rst), .Q(
        \reg_mem[29][29] ) );
  CFD2QXL \reg_mem_reg[29][31]  ( .D(n416), .CP(clk), .CD(rst), .Q(
        \reg_mem[29][31] ) );
  CFD2QXL \reg_mem_reg[31][20]  ( .D(n363), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][20] ) );
  CFD2QXL \reg_mem_reg[31][23]  ( .D(n360), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][23] ) );
  CFD2QXL \reg_mem_reg[31][29]  ( .D(n354), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][29] ) );
  CFD2QXL \reg_mem_reg[31][31]  ( .D(n352), .CP(clk), .CD(rst), .Q(
        \reg_mem[31][31] ) );
  CFD2QXL \reg_mem_reg[30][20]  ( .D(n395), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][20] ) );
  CFD2QXL \reg_mem_reg[30][23]  ( .D(n392), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][23] ) );
  CFD2QXL \reg_mem_reg[30][29]  ( .D(n386), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][29] ) );
  CFD2QXL \reg_mem_reg[30][31]  ( .D(n384), .CP(clk), .CD(rst), .Q(
        \reg_mem[30][31] ) );
  CFD2QXL \reg_mem_reg[9][20]  ( .D(n1067), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][20] ) );
  CFD2QXL \reg_mem_reg[9][23]  ( .D(n1064), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][23] ) );
  CFD2QXL \reg_mem_reg[8][20]  ( .D(n1099), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][20] ) );
  CFD2QXL \reg_mem_reg[8][23]  ( .D(n1096), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][23] ) );
  CFD2QXL \reg_mem_reg[5][20]  ( .D(n1195), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][20] ) );
  CFD2QXL \reg_mem_reg[5][23]  ( .D(n1192), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][23] ) );
  CFD2QXL \reg_mem_reg[5][29]  ( .D(n1186), .CP(clk), .CD(rst), .Q(
        \reg_mem[5][29] ) );
  CFD2QXL \reg_mem_reg[4][20]  ( .D(n1227), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][20] ) );
  CFD2QXL \reg_mem_reg[4][23]  ( .D(n1224), .CP(clk), .CD(rst), .Q(
        \reg_mem[4][23] ) );
  CFD2QXL \reg_mem_reg[3][20]  ( .D(n1259), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][20] ) );
  CFD2QXL \reg_mem_reg[3][23]  ( .D(n1256), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][23] ) );
  CFD2QXL \reg_mem_reg[3][29]  ( .D(n1250), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][29] ) );
  CFD2QXL \reg_mem_reg[3][31]  ( .D(n1248), .CP(clk), .CD(rst), .Q(
        \reg_mem[3][31] ) );
  CFD2QXL \reg_mem_reg[2][15]  ( .D(n1296), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][15] ) );
  CFD2QXL \reg_mem_reg[2][20]  ( .D(n1291), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][20] ) );
  CFD2QXL \reg_mem_reg[2][21]  ( .D(n1290), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][21] ) );
  CFD2QXL \reg_mem_reg[2][23]  ( .D(n1288), .CP(clk), .CD(rst), .Q(
        \reg_mem[2][23] ) );
  CFD2QXL \reg_mem_reg[7][20]  ( .D(n1131), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][20] ) );
  CFD2QXL \reg_mem_reg[7][23]  ( .D(n1128), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][23] ) );
  CFD2QXL \reg_mem_reg[7][29]  ( .D(n1122), .CP(clk), .CD(rst), .Q(
        \reg_mem[7][29] ) );
  CFD2QXL \reg_mem_reg[6][20]  ( .D(n1163), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][20] ) );
  CFD2QXL \reg_mem_reg[6][23]  ( .D(n1160), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][23] ) );
  CFD2QXL \reg_mem_reg[6][29]  ( .D(n1154), .CP(clk), .CD(rst), .Q(
        \reg_mem[6][29] ) );
  CFD2QXL \reg_mem_reg[9][29]  ( .D(n1058), .CP(clk), .CD(rst), .Q(
        \reg_mem[9][29] ) );
  CFD2QXL \reg_mem_reg[1][20]  ( .D(n1323), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][20] ) );
  CFD2QXL \reg_mem_reg[1][23]  ( .D(n1320), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][23] ) );
  CFD2QXL \reg_mem_reg[1][29]  ( .D(n1314), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][29] ) );
  CFD2QXL \reg_mem_reg[1][31]  ( .D(n1312), .CP(clk), .CD(rst), .Q(
        \reg_mem[1][31] ) );
  CFD2QXL \reg_mem_reg[8][29]  ( .D(n1090), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][29] ) );
  CFD2QXL \reg_mem_reg[8][31]  ( .D(n1088), .CP(clk), .CD(rst), .Q(
        \reg_mem[8][31] ) );
  CFD2QXL \reg_mem_reg[0][15]  ( .D(n1360), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][15] ) );
  CFD2QXL \reg_mem_reg[0][20]  ( .D(n1355), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][20] ) );
  CFD2QXL \reg_mem_reg[0][21]  ( .D(n1354), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][21] ) );
  CFD2QXL \reg_mem_reg[0][23]  ( .D(n1352), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][23] ) );
  CFD2QXL \reg_mem_reg[0][29]  ( .D(n1346), .CP(clk), .CD(rst), .Q(
        \reg_mem[0][29] ) );
  CFD1QXL \reg_mem_reg[24][25]  ( .D(n582), .CP(clk), .Q(\reg_mem[24][25] ) );
  CFD2QXL r_type_reg ( .D(net76653), .CP(clk), .CD(rst), .Q(r_type) );
  CFD1QXL \reg_mem_reg[10][26]  ( .D(n1029), .CP(clk), .Q(\reg_mem[10][26] )
         );
  CFD2QXL \prog_count_reg[3]  ( .D(prog_count_c[3]), .CP(clk), .CD(rst), .Q(
        prog_count_o[3]) );
  CFD2QXL i_type_reg ( .D(n5242), .CP(clk), .CD(rst), .Q(i_type) );
  CFD2QXL \regb_addr_reg[3]  ( .D(net82869), .CP(clk), .CD(rst), .Q(
        regb_addr[3]) );
  CFD2QXL \regb_addr_reg[1]  ( .D(net87639), .CP(clk), .CD(rst), .Q(
        regb_addr[1]) );
  CFD2QXL \prog_count_ex_reg[7]  ( .D(n1879), .CP(clk), .CD(rst), .Q(
        prog_count_ex[7]) );
  CFD2QXL \regb_addr_reg[4]  ( .D(net86657), .CP(clk), .CD(rst), .Q(
        regb_addr[4]) );
  CFD2QXL \regb_addr_reg[2]  ( .D(net87720), .CP(clk), .CD(rst), .Q(
        regb_addr[2]) );
  CFD2QXL \regB_reg[30]  ( .D(N202), .CP(clk), .CD(rst), .Q(regB[30]) );
  CFD2QXL \prog_count_reg[4]  ( .D(n1881), .CP(clk), .CD(rst), .Q(
        prog_count_o[4]) );
  CFD2QXL \prog_count_ex_reg[0]  ( .D(n1883), .CP(clk), .CD(rst), .Q(N128) );
  CFD2XL \immi_val_reg[27]  ( .D(n5237), .CP(clk), .CD(rst), .Q(immi_val[27]), 
        .QN(\dp_cluster_0/N36 ) );
  CFD2QXL \prog_count_ex_reg[4]  ( .D(n1886), .CP(clk), .CD(rst), .Q(
        prog_count_ex[4]) );
  CFD2QXL \opcode_ex_reg[3]  ( .D(inst_fetch[3]), .CP(clk), .CD(rst), .Q(
        opcode_ex[3]) );
  CFD2QXL \prog_count_ex_reg[5]  ( .D(n1889), .CP(clk), .CD(rst), .Q(
        prog_count_ex[5]) );
  CFD2QXL \opcode_ex_reg[5]  ( .D(net87691), .CP(clk), .CD(rst), .Q(
        opcode_ex[5]) );
  CFD2QXL \opcode_ex_reg[2]  ( .D(net88116), .CP(clk), .CD(rst), .Q(
        opcode_ex[2]) );
  CFD2QXL j_type_reg ( .D(j_type_c), .CP(clk), .CD(rst), .Q(j_type) );
  CFD2QXL \regc_addr_reg[4]  ( .D(regc_addr_c[4]), .CP(clk), .CD(rst), .Q(
        regc_addr[4]) );
  CFD2QXL \regc_addr_reg[3]  ( .D(regc_addr_c[3]), .CP(clk), .CD(rst), .Q(
        regc_addr[3]) );
  CFD2QXL \regc_addr_reg[2]  ( .D(regc_addr_c[2]), .CP(clk), .CD(rst), .Q(
        regc_addr[2]) );
  CFD2QXL \regc_addr_reg[1]  ( .D(regc_addr_c[1]), .CP(clk), .CD(rst), .Q(
        regc_addr[1]) );
  CFD2QXL \regc_addr_reg[0]  ( .D(regc_addr_c[0]), .CP(clk), .CD(rst), .Q(
        regc_addr[0]) );
  CFD2QXL \opcode_ex_reg[4]  ( .D(inst_fetch[4]), .CP(clk), .CD(rst), .Q(
        opcode_ex[4]) );
  CFD2QX1 \prog_count_ex_reg[1]  ( .D(n1891), .CP(clk), .CD(rst), .Q(N129) );
  CFD2QXL \regB_reg[29]  ( .D(N203), .CP(clk), .CD(rst), .Q(regB[29]) );
  CFD2QX2 \regA_reg[21]  ( .D(N290), .CP(clk), .CD(rst), .Q(regA[21]) );
  CFD1QXL \reg_mem_reg[11][1]  ( .D(n1022), .CP(clk), .Q(\reg_mem[11][1] ) );
  CFD1QXL \reg_mem_reg[15][1]  ( .D(n894), .CP(clk), .Q(\reg_mem[15][1] ) );
  CFD2QXL j_type_wb_reg ( .D(n1896), .CP(clk), .CD(rst), .Q(j_type_wb) );
  CFD2QXL \immi_val_reg[31]  ( .D(n5237), .CP(clk), .CD(rst), .Q(immi_val[31])
         );
  CFD2XL \regA_reg[18]  ( .D(N287), .CP(clk), .CD(rst), .Q(n2125), .QN(n2124)
         );
  CFD2QX1 \immi_val_reg[10]  ( .D(immi_val_c[10]), .CP(clk), .CD(rst), .Q(
        n2118) );
  CFD2QX1 i_type_wb_reg ( .D(i_type_wb_c), .CP(clk), .CD(rst), .Q(i_type_wb)
         );
  CFD2QX1 data_mem_rd_d_reg ( .D(data_mem_rd_o), .CP(clk), .CD(rst), .Q(
        data_mem_rd_d) );
  CFD2XL \regA_reg[1]  ( .D(N270), .CP(clk), .CD(rst), .Q(n2108), .QN(n2107)
         );
  CFD2QXL \regc_addr_mem_reg[4]  ( .D(n1898), .CP(clk), .CD(rst), .Q(
        regc_addr_mem[4]) );
  CFD2QXL \regc_addr_mem_reg[3]  ( .D(n1901), .CP(clk), .CD(rst), .Q(
        regc_addr_mem[3]) );
  CFD2QXL \regc_addr_mem_reg[2]  ( .D(n1904), .CP(clk), .CD(rst), .Q(
        regc_addr_mem[2]) );
  CFD2QXL \regc_addr_mem_reg[1]  ( .D(n1907), .CP(clk), .CD(rst), .Q(
        regc_addr_mem[1]) );
  CFD2QXL \regc_addr_mem_reg[0]  ( .D(n1910), .CP(clk), .CD(rst), .Q(
        regc_addr_mem[0]) );
  CFD2QXL \regb_addr_mem_reg[4]  ( .D(n1913), .CP(clk), .CD(rst), .Q(
        regb_addr_mem[4]) );
  CFD2QXL \regb_addr_mem_reg[3]  ( .D(n1915), .CP(clk), .CD(rst), .Q(
        regb_addr_mem[3]) );
  CFD2QXL \regb_addr_mem_reg[2]  ( .D(n1917), .CP(clk), .CD(rst), .Q(
        regb_addr_mem[2]) );
  CFD2QXL \regb_addr_mem_reg[1]  ( .D(n1919), .CP(clk), .CD(rst), .Q(
        regb_addr_mem[1]) );
  CFD2QXL \regb_addr_mem_reg[0]  ( .D(n1920), .CP(clk), .CD(rst), .Q(
        regb_addr_mem[0]) );
  CFD2QXL \prog_count_de_reg[0]  ( .D(n1922), .CP(clk), .CD(rst), .Q(
        prog_count_de[0]) );
  CFD2QXL \prog_count_de_reg[7]  ( .D(n1924), .CP(clk), .CD(rst), .Q(
        prog_count_de[7]) );
  CFD2QXL \prog_count_de_reg[4]  ( .D(n1927), .CP(clk), .CD(rst), .Q(
        prog_count_de[4]) );
  CFD2QXL \prog_count_de_reg[5]  ( .D(n1929), .CP(clk), .CD(rst), .Q(
        prog_count_de[5]) );
  CFD2QXL \prog_count_de_reg[6]  ( .D(n1930), .CP(clk), .CD(rst), .Q(
        prog_count_de[6]) );
  CFD2QXL r_type_mem_reg ( .D(n1931), .CP(clk), .CD(rst), .Q(r_type_mem) );
  CFD2QXL \prog_count_de_reg[1]  ( .D(n1932), .CP(clk), .CD(rst), .Q(
        prog_count_de[1]) );
  CFD2QXL \prog_count_de_reg[2]  ( .D(n1934), .CP(clk), .CD(rst), .Q(
        prog_count_de[2]) );
  CFD2QXL \prog_count_de_reg[3]  ( .D(n1935), .CP(clk), .CD(rst), .Q(
        prog_count_de[3]) );
  CFD2QX2 \regB_reg[12]  ( .D(N220), .CP(clk), .CD(rst), .Q(regB[12]) );
  CFD2QX2 \regB_reg[8]  ( .D(N224), .CP(clk), .CD(rst), .Q(regB[8]) );
  CFD2QX2 \regB_reg[21]  ( .D(N211), .CP(clk), .CD(rst), .Q(regB[21]) );
  CFD2QX2 \regB_reg[25]  ( .D(N207), .CP(clk), .CD(rst), .Q(regB[25]) );
  CFD2QX2 \regB_reg[10]  ( .D(N222), .CP(clk), .CD(rst), .Q(regB[10]) );
  CFD2QX2 \regB_reg[7]  ( .D(N225), .CP(clk), .CD(rst), .Q(regB[7]) );
  CFD2QX2 \regB_reg[0]  ( .D(N232), .CP(clk), .CD(rst), .Q(regB[0]) );
  CFD2QX2 \regB_reg[20]  ( .D(N212), .CP(clk), .CD(rst), .Q(regB[20]) );
  CFD2QX2 \regB_reg[19]  ( .D(N213), .CP(clk), .CD(rst), .Q(regB[19]) );
  CFD2QX2 \regB_reg[22]  ( .D(N210), .CP(clk), .CD(rst), .Q(regB[22]) );
  CFD2QX2 \regB_reg[15]  ( .D(N217), .CP(clk), .CD(rst), .Q(regB[15]) );
  CFD2QX2 \regB_reg[26]  ( .D(N206), .CP(clk), .CD(rst), .Q(regB[26]) );
  CFD2QX1 \immi_val_reg[4]  ( .D(immi_val_c[4]), .CP(clk), .CD(rst), .Q(n2061)
         );
  CFD2XL \regA_reg[24]  ( .D(N293), .CP(clk), .CD(rst), .Q(n2057), .QN(n2056)
         );
  CFD2QX2 \regB_reg[28]  ( .D(N204), .CP(clk), .CD(rst), .Q(regB[28]) );
  CFD2QX2 \regB_reg[24]  ( .D(N208), .CP(clk), .CD(rst), .Q(regB[24]) );
  CFD2X2 \regB_reg[17]  ( .D(N215), .CP(clk), .CD(rst), .Q(n2051) );
  CFD2X2 \regB_reg[5]  ( .D(N227), .CP(clk), .CD(rst), .Q(n2049), .QN(n2048)
         );
  CFD2X1 \regA_reg[29]  ( .D(N298), .CP(clk), .CD(rst), .Q(n2029) );
  CFD2QX2 \regB_reg[6]  ( .D(N226), .CP(clk), .CD(rst), .Q(regB[6]) );
  CFD2X2 \regA_reg[17]  ( .D(N286), .CP(clk), .CD(rst), .Q(n2024), .QN(n2023)
         );
  CFD2XL \regB_reg[23]  ( .D(N209), .CP(clk), .CD(rst), .Q(n2020), .QN(n2019)
         );
  CAOR2X1 U833 ( .A(\reg_mem[19][4] ), .B(n214), .C(net81907), .D(net83073), 
        .Z(n763) );
  CAOR2X1 U865 ( .A(\reg_mem[18][4] ), .B(n1507), .C(net81947), .D(net83072), 
        .Z(n795) );
  CAOR2X1 U897 ( .A(\reg_mem[17][4] ), .B(n1505), .C(net81987), .D(n186), .Z(
        n827) );
  CAOR2X1 U929 ( .A(\reg_mem[16][4] ), .B(n1509), .C(net82027), .D(net83073), 
        .Z(n859) );
  CAOR2X1 U835 ( .A(\reg_mem[19][2] ), .B(n214), .C(net81905), .D(net83077), 
        .Z(n765) );
  CAOR2X1 U867 ( .A(\reg_mem[18][2] ), .B(n1507), .C(net81945), .D(net83076), 
        .Z(n797) );
  CAOR2X1 U899 ( .A(\reg_mem[17][2] ), .B(n1505), .C(net81985), .D(n188), .Z(
        n829) );
  CAOR2X1 U931 ( .A(\reg_mem[16][2] ), .B(n1509), .C(net82025), .D(net83077), 
        .Z(n861) );
  CAOR2X1 U1242 ( .A(\reg_mem[6][11] ), .B(n232), .C(net82425), .D(net83058), 
        .Z(n1172) );
  CAOR2X1 U1210 ( .A(\reg_mem[7][11] ), .B(net82377), .C(net82385), .D(
        net83059), .Z(n1140) );
  CAOR2X1 U1274 ( .A(\reg_mem[5][11] ), .B(net82457), .C(net82473), .D(n179), 
        .Z(n1204) );
  CAOR2X1 U1306 ( .A(\reg_mem[4][11] ), .B(net82497), .C(net82513), .D(
        net83059), .Z(n1236) );
  CAOR2X1 U1336 ( .A(\reg_mem[3][13] ), .B(net82539), .C(net82549), .D(
        net83054), .Z(n1266) );
  CAOR2X1 U1368 ( .A(\reg_mem[2][13] ), .B(net82579), .C(net82591), .D(n177), 
        .Z(n1298) );
  CAOR2X1 U1400 ( .A(\reg_mem[1][13] ), .B(net82619), .C(net82625), .D(
        net83055), .Z(n1330) );
  CAOR2X1 U1450 ( .A(\reg_mem[0][13] ), .B(n1530), .C(net82665), .D(net83054), 
        .Z(n1362) );
  CFD2X2 \regB_reg[4]  ( .D(N228), .CP(clk), .CD(rst), .Q(n2110) );
  CFD2X2 \regB_reg[2]  ( .D(N230), .CP(clk), .CD(rst), .Q(n2047) );
  CFD2X2 \regB_reg[11]  ( .D(N221), .CP(clk), .CD(rst), .Q(n2033) );
  CFD2X2 \regB_reg[13]  ( .D(N219), .CP(clk), .CD(rst), .Q(n2026) );
  CFD1QX1 \reg_mem_reg[20][29]  ( .D(n706), .CP(clk), .Q(\reg_mem[20][29] ) );
  CFD2X1 \regA_reg[8]  ( .D(N277), .CP(clk), .CD(rst), .Q(n2059) );
  CFD2X4 \regA_reg[26]  ( .D(N295), .CP(clk), .CD(rst), .Q(n2015), .QN(n2014)
         );
  CFD2XL \immi_val_reg[25]  ( .D(immi_val_c[25]), .CP(clk), .CD(rst), .Q(
        immi_val[25]), .QN(\dp_cluster_0/N38 ) );
  CFD2XL \immi_val_reg[24]  ( .D(immi_val_c[24]), .CP(clk), .CD(rst), .Q(
        immi_val[24]), .QN(\dp_cluster_0/N39 ) );
  CFD2XL \immi_val_reg[30]  ( .D(n5237), .CP(clk), .CD(rst), .Q(immi_val[30]), 
        .QN(\dp_cluster_0/N33 ) );
  CFD2XL \immi_val_reg[29]  ( .D(n5237), .CP(clk), .CD(rst), .Q(immi_val[29]), 
        .QN(\dp_cluster_0/N34 ) );
  CFD2XL \immi_val_reg[28]  ( .D(n5237), .CP(clk), .CD(rst), .Q(immi_val[28]), 
        .QN(\dp_cluster_0/N35 ) );
  CFD1XL \reg_mem_reg[23][23]  ( .D(n616), .CP(clk), .Q(\reg_mem[23][23] ), 
        .QN(n4791) );
  CFD4XL \reg_mem_reg[29][15]  ( .D(n432), .CP(clk), .SD(rst), .Q(
        \reg_mem[29][15] ), .QN(n4421) );
  CFD4XL \reg_mem_reg[29][14]  ( .D(n433), .CP(clk), .SD(rst), .Q(
        \reg_mem[29][14] ), .QN(n4359) );
  CFD4XL \reg_mem_reg[29][13]  ( .D(n434), .CP(clk), .SD(rst), .Q(
        \reg_mem[29][13] ), .QN(n4317) );
  CFD4XL \reg_mem_reg[29][12]  ( .D(n435), .CP(clk), .SD(rst), .Q(
        \reg_mem[29][12] ), .QN(n4283) );
  CFD4XL \reg_mem_reg[29][11]  ( .D(n436), .CP(clk), .SD(rst), .Q(
        \reg_mem[29][11] ), .QN(n4241) );
  CFD4XL \reg_mem_reg[29][10]  ( .D(n437), .CP(clk), .SD(rst), .Q(
        \reg_mem[29][10] ), .QN(n4207) );
  CFD4XL \reg_mem_reg[29][9]  ( .D(n438), .CP(clk), .SD(rst), .Q(
        \reg_mem[29][9] ), .QN(n4163) );
  CFD4XL \reg_mem_reg[29][8]  ( .D(n439), .CP(clk), .SD(rst), .Q(
        \reg_mem[29][8] ), .QN(n4119) );
  CFD4XL \reg_mem_reg[29][7]  ( .D(n440), .CP(clk), .SD(rst), .Q(
        \reg_mem[29][7] ), .QN(n4073) );
  CFD4XL \reg_mem_reg[29][6]  ( .D(n441), .CP(clk), .SD(rst), .Q(
        \reg_mem[29][6] ), .QN(n4029) );
  CFD4XL \reg_mem_reg[29][5]  ( .D(n442), .CP(clk), .SD(rst), .Q(
        \reg_mem[29][5] ), .QN(n3985) );
  CFD4XL \reg_mem_reg[29][4]  ( .D(n443), .CP(clk), .SD(rst), .Q(
        \reg_mem[29][4] ), .QN(n3945) );
  CFD4XL \reg_mem_reg[29][3]  ( .D(n444), .CP(clk), .SD(rst), .Q(
        \reg_mem[29][3] ), .QN(n3909) );
  CFD4XL \reg_mem_reg[29][2]  ( .D(n445), .CP(clk), .SD(rst), .Q(
        \reg_mem[29][2] ), .QN(n3869) );
  CFD4XL \reg_mem_reg[29][1]  ( .D(n446), .CP(clk), .SD(rst), .Q(
        \reg_mem[29][1] ), .QN(n3833) );
  CFD4XL \reg_mem_reg[29][0]  ( .D(n447), .CP(clk), .SD(rst), .Q(
        \reg_mem[29][0] ), .QN(n3789) );
  CFD4XL \reg_mem_reg[31][7]  ( .D(n376), .CP(clk), .SD(rst), .Q(
        \reg_mem[31][7] ), .QN(n4075) );
  CFD4XL \reg_mem_reg[31][5]  ( .D(n378), .CP(clk), .SD(rst), .Q(
        \reg_mem[31][5] ), .QN(n3987) );
  CFD4XL \reg_mem_reg[4][2]  ( .D(n1245), .CP(clk), .SD(rst), .Q(
        \reg_mem[4][2] ) );
  CFD4XL \reg_mem_reg[4][1]  ( .D(n1246), .CP(clk), .SD(rst), .Q(
        \reg_mem[4][1] ) );
  CFD2XL \prog_count_reg[2]  ( .D(n1467), .CP(clk), .CD(rst), .Q(
        prog_count_o[2]), .QN(n3480) );
  CFD2X2 \regB_reg[3]  ( .D(N229), .CP(clk), .CD(rst), .Q(n1685), .QN(n1684)
         );
  CFD2X1 \regA_reg[25]  ( .D(N294), .CP(clk), .CD(rst), .Q(n2036), .QN(n2035)
         );
  CFD2QX2 \regB_reg[18]  ( .D(N214), .CP(clk), .CD(rst), .Q(regB[18]) );
  CFD2QX2 \regB_reg[14]  ( .D(N218), .CP(clk), .CD(rst), .Q(regB[14]) );
  CFD2X1 \immi_val_reg[18]  ( .D(immi_val_c[18]), .CP(clk), .CD(rst), .Q(
        immi_val[18]), .QN(\dp_cluster_0/N45 ) );
  CFD2QX1 \prog_count_ex_reg[2]  ( .D(n1689), .CP(clk), .CD(rst), .Q(
        prog_count_ex[2]) );
  CFD2QX1 \prog_count_ex_reg[3]  ( .D(n1687), .CP(clk), .CD(rst), .Q(
        prog_count_ex[3]) );
  CFD2QX1 \regA_reg[13]  ( .D(N282), .CP(clk), .CD(rst), .Q(regA[13]) );
  CFD2QX1 \regB_reg[31]  ( .D(N201), .CP(clk), .CD(rst), .Q(regB[31]) );
  CFD2QX1 \regB_reg[9]  ( .D(N223), .CP(clk), .CD(rst), .Q(regB[9]) );
  CFD2X1 \regB_reg[16]  ( .D(N216), .CP(clk), .CD(rst), .Q(n2106) );
  CFD1QXL \reg_mem_reg[26][26]  ( .D(n1937), .CP(clk), .Q(\reg_mem[26][26] )
         );
  CFD2QX1 \prog_count_ex_reg[6]  ( .D(n1894), .CP(clk), .CD(rst), .Q(
        prog_count_ex[6]) );
  CFD4XL \reg_mem_reg[4][0]  ( .D(n1247), .CP(clk), .SD(rst), .Q(
        \reg_mem[4][0] ), .QN(n1594) );
  CFD2QX2 \regA_reg[4]  ( .D(N273), .CP(clk), .CD(rst), .Q(regA[4]) );
  CFD2X2 \regA_reg[14]  ( .D(N283), .CP(clk), .CD(rst), .Q(n1494), .QN(n1493)
         );
  CFD2X2 \regA_reg[12]  ( .D(N281), .CP(clk), .CD(rst), .Q(n1475), .QN(n1474)
         );
  CFD2QX1 \regA_reg[27]  ( .D(N296), .CP(clk), .CD(rst), .Q(regA[27]) );
  CFD2QX1 \regA_reg[15]  ( .D(N284), .CP(clk), .CD(rst), .Q(regA[15]) );
  CFD2QX2 \regB_reg[27]  ( .D(N205), .CP(clk), .CD(rst), .Q(regB[27]) );
  CFD2QX1 \regB_reg[1]  ( .D(N231), .CP(clk), .CD(rst), .Q(regB[1]) );
  CFD2X2 \regA_reg[0]  ( .D(N269), .CP(clk), .CD(rst), .Q(n1387), .QN(n1386)
         );
  CFD2X2 \regA_reg[20]  ( .D(N289), .CP(clk), .CD(rst), .Q(n1379), .QN(n1378)
         );
  CMXI2X1 U1524 ( .A0(n2965), .A1(n2966), .S(n1470), .Z(n2970) );
  CMXI2X1 U1525 ( .A0(n3550), .A1(n3549), .S(n2191), .Z(n3551) );
  CIVX2 U1526 ( .A(n1378), .Z(n1380) );
  CMXI2X1 U1527 ( .A0(n3247), .A1(n3246), .S(n2097), .Z(n3249) );
  CNR2IX1 U1528 ( .B(n3615), .A(n2778), .Z(n2784) );
  CMXI2X1 U1529 ( .A0(n3472), .A1(n3473), .S(n3615), .Z(N273) );
  CMXI2X1 U1530 ( .A0(n3471), .A1(n3470), .S(n1390), .Z(n3473) );
  CNIVX3 U1531 ( .A(net87511), .Z(net87525) );
  CAN2XL U1532 ( .A(n2886), .B(n2176), .Z(n1669) );
  CMXI2X1 U1533 ( .A0(\reg_mem[20][18] ), .A1(\reg_mem[4][18] ), .S(n1382), 
        .Z(n2948) );
  CIVX2 U1534 ( .A(n2086), .Z(n1382) );
  CNIVX3 U1535 ( .A(n2076), .Z(n2081) );
  CNIVX2 U1536 ( .A(net87380), .Z(net87411) );
  CMXI2XL U1537 ( .A0(\reg_mem[5][27] ), .A1(\reg_mem[21][27] ), .S(n2103), 
        .Z(n2614) );
  CMXI2XL U1538 ( .A0(n4394), .A1(n4424), .S(n2103), .Z(n3059) );
  CMXI2XL U1539 ( .A0(\reg_mem[11][31] ), .A1(\reg_mem[27][31] ), .S(n2103), 
        .Z(n3650) );
  CMXI2XL U1540 ( .A0(\reg_mem[3][31] ), .A1(\reg_mem[19][31] ), .S(n2103), 
        .Z(n3668) );
  CMXI2XL U1541 ( .A0(n4937), .A1(n4967), .S(n2103), .Z(n2633) );
  CMXI2XL U1542 ( .A0(\reg_mem[0][30] ), .A1(\reg_mem[16][30] ), .S(n2103), 
        .Z(n3606) );
  CMXI2X1 U1543 ( .A0(\reg_mem[16][20] ), .A1(\reg_mem[24][20] ), .S(net87522), 
        .Z(n2885) );
  CNIVX2 U1544 ( .A(net87234), .Z(n1381) );
  CMXI2XL U1545 ( .A0(n2985), .A1(n2986), .S(n2164), .Z(n2987) );
  CIVX2 U1546 ( .A(n2086), .Z(n2072) );
  CMXI2XL U1547 ( .A0(n2971), .A1(n2972), .S(n1531), .Z(n1983) );
  CNIVX3 U1548 ( .A(net87380), .Z(net87412) );
  CNIVX2 U1549 ( .A(net87234), .Z(net87242) );
  CMXI2XL U1550 ( .A0(n3410), .A1(n3409), .S(n1389), .Z(n3426) );
  CNIVX3 U1551 ( .A(net87514), .Z(net87523) );
  CIVX1 U1552 ( .A(n2172), .Z(n1383) );
  CIVX3 U1553 ( .A(n2167), .Z(n2172) );
  CND2X1 U1554 ( .A(n2887), .B(n2133), .Z(n2134) );
  CMXI2XL U1555 ( .A0(n2958), .A1(n2957), .S(n1389), .Z(n1984) );
  CIVX3 U1556 ( .A(n1381), .Z(n1384) );
  CIVX4 U1557 ( .A(n1384), .Z(n1385) );
  CNIVX2 U1558 ( .A(net87242), .Z(net87267) );
  CMXI2XL U1559 ( .A0(\reg_mem[8][1] ), .A1(\reg_mem[12][1] ), .S(net87243), 
        .Z(n3575) );
  CANR2X1 U1560 ( .A(N198), .B(n2140), .C(n1533), .D(n2545), .Z(n2542) );
  CIVDX1 U1561 ( .A(net87540), .Z0(net87508), .Z1(n1389) );
  CIVX4 U1562 ( .A(n1386), .Z(n1388) );
  CND2IX1 U1563 ( .B(n3811), .A(net87243), .Z(n2131) );
  CNIVX3 U1564 ( .A(net87512), .Z(net87533) );
  CNIVX3 U1565 ( .A(net87514), .Z(net87532) );
  CNIVX4 U1566 ( .A(net87516), .Z(net87541) );
  CIVX2 U1567 ( .A(n1458), .Z(n1390) );
  CNR2IX2 U1568 ( .B(n2820), .A(n2819), .Z(n2821) );
  CMXI2XL U1569 ( .A0(n3553), .A1(n3554), .S(net87508), .Z(n3555) );
  CMXI2XL U1570 ( .A0(n2991), .A1(n2992), .S(n2039), .Z(n2996) );
  CMXI2X1 U1571 ( .A0(\reg_mem[19][20] ), .A1(\reg_mem[27][20] ), .S(net87533), 
        .Z(n2889) );
  CMXI2X1 U1572 ( .A0(n2890), .A1(n2889), .S(n2182), .Z(n2894) );
  CMXI2X1 U1573 ( .A0(n2995), .A1(n2996), .S(n1392), .Z(n3004) );
  CNIVX1 U1574 ( .A(net87238), .Z(net87262) );
  CNIVX1 U1575 ( .A(net87241), .Z(net87278) );
  CNIVX2 U1576 ( .A(net87513), .Z(net87520) );
  CNIVX2 U1577 ( .A(net87513), .Z(net87538) );
  CIVX2 U1578 ( .A(n1392), .Z(n1391) );
  CIVX3 U1579 ( .A(net87279), .Z(n1392) );
  CND3X1 U1580 ( .A(n3674), .B(n3673), .C(n3672), .Z(n3684) );
  CND2IX1 U1581 ( .B(n2543), .A(n2542), .Z(N298) );
  CNR2IX1 U1582 ( .B(n3615), .A(n2537), .Z(n2543) );
  CMXI2X1 U1583 ( .A0(n2064), .A1(n2063), .S(n1458), .Z(n2151) );
  CMXI2X1 U1584 ( .A0(n2517), .A1(n2518), .S(n1392), .Z(n2519) );
  CMXI2XL U1585 ( .A0(net79033), .A1(net79032), .S(n2175), .Z(n3546) );
  CIVX3 U1586 ( .A(n2175), .Z(n2183) );
  CNIVX3 U1587 ( .A(n2076), .Z(n2098) );
  CANR2XL U1588 ( .A(alu_op_c[6]), .B(n3750), .C(regA[6]), .D(n3739), .Z(n3346) );
  CIVXL U1589 ( .A(alu_op_c[6]), .Z(n3379) );
  CNIVXL U1590 ( .A(regB[30]), .Z(n1699) );
  CND2IXL U1591 ( .B(n3612), .A(n3611), .Z(n3613) );
  CMXI2XL U1592 ( .A0(n4663), .A1(n4693), .S(n2080), .Z(n2835) );
  CMXI2X1 U1593 ( .A0(n5213), .A1(n5214), .S(net87990), .Z(N201) );
  CMXI2XL U1594 ( .A0(n4538), .A1(n4537), .S(net87626), .Z(n4544) );
  CMXI2XL U1595 ( .A0(n1393), .A1(n1394), .S(net87790), .Z(net77967) );
  CIVX20 U1596 ( .A(\reg_mem[4][13] ), .Z(n1393) );
  CIVX20 U1597 ( .A(\reg_mem[5][13] ), .Z(n1394) );
  CMXI2XL U1598 ( .A0(n1395), .A1(n1396), .S(net87790), .Z(n4300) );
  CIVX20 U1599 ( .A(\reg_mem[12][13] ), .Z(n1395) );
  CIVX20 U1600 ( .A(\reg_mem[13][13] ), .Z(n1396) );
  CMXI2XL U1601 ( .A0(n1397), .A1(n1398), .S(net87797), .Z(n5133) );
  CIVX20 U1602 ( .A(\reg_mem[18][30] ), .Z(n1397) );
  CIVX20 U1603 ( .A(\reg_mem[19][30] ), .Z(n1398) );
  CMXI2XL U1604 ( .A0(n4260), .A1(n4259), .S(net87629), .Z(n4266) );
  CMXI2XL U1605 ( .A0(n1399), .A1(n1400), .S(net87798), .Z(n4049) );
  CIVX20 U1606 ( .A(\reg_mem[10][7] ), .Z(n1399) );
  CIVX20 U1607 ( .A(\reg_mem[11][7] ), .Z(n1400) );
  CMXI2XL U1608 ( .A0(n1401), .A1(n1402), .S(net87790), .Z(n4092) );
  CIVX20 U1609 ( .A(\reg_mem[4][8] ), .Z(n1401) );
  CIVX20 U1610 ( .A(\reg_mem[5][8] ), .Z(n1402) );
  CMXI2XL U1611 ( .A0(n1403), .A1(n1404), .S(net87790), .Z(n4524) );
  CIVX20 U1612 ( .A(\reg_mem[4][18] ), .Z(n1403) );
  CIVX20 U1613 ( .A(\reg_mem[5][18] ), .Z(n1404) );
  CMXI2XL U1614 ( .A0(n1405), .A1(n1406), .S(net87802), .Z(n4020) );
  CIVX20 U1615 ( .A(\reg_mem[20][6] ), .Z(n1405) );
  CIVX20 U1616 ( .A(\reg_mem[21][6] ), .Z(n1406) );
  CNIVXL U1617 ( .A(prog_count_c[2]), .Z(n1467) );
  CMXI2XL U1618 ( .A0(n5021), .A1(n5022), .S(n1453), .Z(N205) );
  CMXI2XL U1619 ( .A0(n1407), .A1(n1408), .S(net87800), .Z(n3810) );
  CIVX20 U1620 ( .A(\reg_mem[8][1] ), .Z(n1407) );
  CIVX20 U1621 ( .A(\reg_mem[9][1] ), .Z(n1408) );
  CMXI2XL U1622 ( .A0(n4528), .A1(n4527), .S(net87623), .Z(n4534) );
  CIVXL U1623 ( .A(immi_val[2]), .Z(n1409) );
  CMXI2XL U1624 ( .A0(n2489), .A1(n2488), .S(n1532), .Z(n2490) );
  CMXI2XL U1625 ( .A0(n2481), .A1(n2480), .S(n1385), .Z(n2489) );
  CMXI2XL U1626 ( .A0(n2505), .A1(n2506), .S(n3615), .Z(N269) );
  CMXI2XL U1627 ( .A0(n2491), .A1(n2490), .S(n2092), .Z(n2506) );
  CMXI2XL U1628 ( .A0(n1410), .A1(n1411), .S(net87804), .Z(n3775) );
  CIVX20 U1629 ( .A(\reg_mem[18][0] ), .Z(n1410) );
  CIVX20 U1630 ( .A(\reg_mem[19][0] ), .Z(n1411) );
  CMXI2XL U1631 ( .A0(n1412), .A1(n1413), .S(net87797), .Z(n4345) );
  CIVX20 U1632 ( .A(\reg_mem[18][14] ), .Z(n1412) );
  CIVX20 U1633 ( .A(\reg_mem[19][14] ), .Z(n1413) );
  CMXI2XL U1634 ( .A0(n1414), .A1(n1415), .S(net87793), .Z(n4228) );
  CIVX20 U1635 ( .A(\reg_mem[16][11] ), .Z(n1414) );
  CIVX20 U1636 ( .A(\reg_mem[17][11] ), .Z(n1415) );
  CMXI2XL U1637 ( .A0(n1416), .A1(n1417), .S(net87807), .Z(n4626) );
  CIVX20 U1638 ( .A(\reg_mem[20][20] ), .Z(n1416) );
  CIVX20 U1639 ( .A(\reg_mem[21][20] ), .Z(n1417) );
  CIVX2 U1640 ( .A(n2168), .Z(n2188) );
  CMXI2XL U1641 ( .A0(n4218), .A1(n4217), .S(net86657), .Z(N222) );
  CIVX4 U1642 ( .A(net86657), .Z(n1453) );
  CMXI2XL U1643 ( .A0(n1418), .A1(n1419), .S(net87795), .Z(n4480) );
  CIVX20 U1644 ( .A(\reg_mem[4][17] ), .Z(n1418) );
  CIVX20 U1645 ( .A(\reg_mem[5][17] ), .Z(n1419) );
  CMXI2XL U1646 ( .A0(n1420), .A1(n1421), .S(net87800), .Z(n4622) );
  CIVX20 U1647 ( .A(\reg_mem[16][20] ), .Z(n1420) );
  CIVX20 U1648 ( .A(\reg_mem[17][20] ), .Z(n1421) );
  CMXI2XL U1649 ( .A0(n1422), .A1(n1423), .S(net87804), .Z(n4220) );
  CIVX20 U1650 ( .A(\reg_mem[8][11] ), .Z(n1422) );
  CIVX20 U1651 ( .A(\reg_mem[9][11] ), .Z(n1423) );
  CMXI2XL U1652 ( .A0(n1424), .A1(n1425), .S(net87791), .Z(n4224) );
  CIVX20 U1653 ( .A(\reg_mem[12][11] ), .Z(n1424) );
  CIVX20 U1654 ( .A(\reg_mem[13][11] ), .Z(n1425) );
  CMXI2X1 U1655 ( .A0(n4219), .A1(n4220), .S(net88166), .Z(n4226) );
  CIVX3 U1656 ( .A(net87639), .Z(net88166) );
  CMXI2X1 U1657 ( .A0(n4223), .A1(n4224), .S(net88166), .Z(n4225) );
  CMXI2XL U1658 ( .A0(n1426), .A1(n1427), .S(net87799), .Z(n4336) );
  CIVX20 U1659 ( .A(\reg_mem[8][14] ), .Z(n1426) );
  CIVX20 U1660 ( .A(\reg_mem[9][14] ), .Z(n1427) );
  CMXI2X1 U1661 ( .A0(n4335), .A1(n4336), .S(net88166), .Z(n4342) );
  CMXI2XL U1662 ( .A0(n1428), .A1(n1429), .S(net87800), .Z(n4227) );
  CIVX20 U1663 ( .A(\reg_mem[18][11] ), .Z(n1428) );
  CIVX20 U1664 ( .A(\reg_mem[19][11] ), .Z(n1429) );
  CMXI2XL U1665 ( .A0(n1430), .A1(n1431), .S(net87807), .Z(n4616) );
  CIVX20 U1666 ( .A(\reg_mem[12][20] ), .Z(n1430) );
  CIVX20 U1667 ( .A(\reg_mem[13][20] ), .Z(n1431) );
  CMXI2XL U1668 ( .A0(n1432), .A1(n1433), .S(net87791), .Z(n4537) );
  CIVX20 U1669 ( .A(\reg_mem[18][18] ), .Z(n1432) );
  CIVX20 U1670 ( .A(\reg_mem[19][18] ), .Z(n1433) );
  CMXI2XL U1671 ( .A0(n1434), .A1(n1435), .S(net87793), .Z(n4538) );
  CIVX20 U1672 ( .A(\reg_mem[16][18] ), .Z(n1434) );
  CIVX20 U1673 ( .A(\reg_mem[17][18] ), .Z(n1435) );
  CMXI2XL U1674 ( .A0(n3600), .A1(n3599), .S(n2193), .Z(n3601) );
  CND2IXL U1675 ( .B(n3604), .A(n3603), .Z(n3614) );
  CMXI2XL U1676 ( .A0(n3602), .A1(n3601), .S(net87265), .Z(n3603) );
  CND2XL U1677 ( .A(n1988), .B(n1946), .Z(n1943) );
  CMXI2XL U1678 ( .A0(n1436), .A1(n1437), .S(net87799), .Z(n4528) );
  CIVX20 U1679 ( .A(\reg_mem[8][18] ), .Z(n1436) );
  CIVX20 U1680 ( .A(\reg_mem[9][18] ), .Z(n1437) );
  CMXI2XL U1681 ( .A0(n5020), .A1(n5019), .S(net82867), .Z(n5021) );
  CNIVX3 U1682 ( .A(net15031), .Z(net82867) );
  CMXI2X1 U1683 ( .A0(n1438), .A1(n1439), .S(net87795), .Z(n4154) );
  CIVX20 U1684 ( .A(\reg_mem[20][9] ), .Z(n1438) );
  CIVX20 U1685 ( .A(\reg_mem[21][9] ), .Z(n1439) );
  CMXI2XL U1686 ( .A0(n4072), .A1(n4071), .S(net87637), .Z(n4080) );
  CMXI2X1 U1687 ( .A0(n1440), .A1(n1441), .S(net87791), .Z(n4350) );
  CIVX20 U1688 ( .A(\reg_mem[20][14] ), .Z(n1440) );
  CIVX20 U1689 ( .A(\reg_mem[21][14] ), .Z(n1441) );
  CMXI2XL U1690 ( .A0(n1442), .A1(n1443), .S(net87790), .Z(n3966) );
  CIVX20 U1691 ( .A(\reg_mem[12][5] ), .Z(n1442) );
  CIVX20 U1692 ( .A(\reg_mem[13][5] ), .Z(n1443) );
  CMXI2XL U1693 ( .A0(n1444), .A1(n1445), .S(net87799), .Z(n4140) );
  CIVX20 U1694 ( .A(\reg_mem[8][9] ), .Z(n1444) );
  CIVX20 U1695 ( .A(\reg_mem[9][9] ), .Z(n1445) );
  CMXI2X1 U1696 ( .A0(n3244), .A1(n3245), .S(n1531), .Z(n3246) );
  CMXI2XL U1697 ( .A0(n1446), .A1(n1447), .S(net87793), .Z(n4144) );
  CIVX20 U1698 ( .A(\reg_mem[12][9] ), .Z(n1446) );
  CIVX20 U1699 ( .A(\reg_mem[13][9] ), .Z(n1447) );
  CMXI2XL U1700 ( .A0(n3960), .A1(n3959), .S(net87723), .Z(n3970) );
  CMXI2X1 U1701 ( .A0(n4143), .A1(n4144), .S(n1988), .Z(n4145) );
  CMXI2XL U1702 ( .A0(n1448), .A1(n1449), .S(net87800), .Z(n4327) );
  CIVX20 U1703 ( .A(\reg_mem[2][14] ), .Z(n1448) );
  CIVX20 U1704 ( .A(\reg_mem[3][14] ), .Z(n1449) );
  CIVX2 U1705 ( .A(n2172), .Z(n1450) );
  CMXI2XL U1706 ( .A0(n1451), .A1(n1452), .S(net87807), .Z(n4346) );
  CIVX20 U1707 ( .A(\reg_mem[16][14] ), .Z(n1451) );
  CIVX20 U1708 ( .A(\reg_mem[17][14] ), .Z(n1452) );
  CIVX8 U1709 ( .A(net87280), .Z(net87233) );
  CNIVX4 U1710 ( .A(net87241), .Z(net87280) );
  CMXI2XL U1711 ( .A0(alu_op_c[13]), .A1(n3144), .S(n1534), .Z(n3145) );
  CMXI2X1 U1712 ( .A0(n4369), .A1(n4370), .S(n1453), .Z(N218) );
  CMXI2X1 U1713 ( .A0(n1454), .A1(n1455), .S(net87793), .Z(n4150) );
  CIVX20 U1714 ( .A(\reg_mem[16][9] ), .Z(n1454) );
  CIVX20 U1715 ( .A(\reg_mem[17][9] ), .Z(n1455) );
  COND3XL U1716 ( .A(n2271), .B(n3184), .C(n3183), .D(n3182), .Z(n3186) );
  CMXI2XL U1717 ( .A0(n2675), .A1(n2674), .S(n2179), .Z(n2676) );
  CNIVX4 U1718 ( .A(n2053), .Z(n1456) );
  CNIVX1 U1719 ( .A(n2053), .Z(n2068) );
  CND2X1 U1720 ( .A(n2632), .B(n2631), .Z(n2668) );
  CMXI2X1 U1721 ( .A0(n3103), .A1(n3104), .S(n1470), .Z(n3105) );
  CMXI2X1 U1722 ( .A0(n5063), .A1(n5064), .S(net87990), .Z(N204) );
  CMXI2X1 U1723 ( .A0(\reg_mem[14][13] ), .A1(\reg_mem[6][13] ), .S(n1531), 
        .Z(n3120) );
  COND3XL U1724 ( .A(n2627), .B(n2626), .C(n2624), .D(n2625), .Z(N296) );
  CMXI2XL U1725 ( .A0(n3584), .A1(n3583), .S(n2185), .Z(n3585) );
  CMXI2XL U1726 ( .A0(n3278), .A1(n3277), .S(net87258), .Z(n3279) );
  CMXI2XL U1727 ( .A0(n3276), .A1(n3275), .S(n2192), .Z(n3277) );
  CMXI2XL U1728 ( .A0(n4292), .A1(n4291), .S(net82863), .Z(n4293) );
  CMX2X1 U1729 ( .A0(n1683), .A1(n1682), .S(n1988), .Z(n4438) );
  CNIVX2 U1730 ( .A(net87241), .Z(net87277) );
  CNIVX2 U1731 ( .A(net87241), .Z(net87281) );
  CNIVX3 U1732 ( .A(net87241), .Z(net87279) );
  CAN2X1 U1733 ( .A(net87233), .B(net87540), .Z(n2148) );
  CMXI2XL U1734 ( .A0(n3108), .A1(n3107), .S(n2201), .Z(n3112) );
  CMXI2XL U1735 ( .A0(\reg_mem[0][16] ), .A1(\reg_mem[8][16] ), .S(net87537), 
        .Z(n3009) );
  CMXI2XL U1736 ( .A0(\reg_mem[5][8] ), .A1(\reg_mem[4][8] ), .S(n2066), .Z(
        n1535) );
  CIVXL U1737 ( .A(n3556), .Z(n1457) );
  CND2XL U1738 ( .A(n3615), .B(n1458), .Z(n1459) );
  CIVXL U1739 ( .A(n2101), .Z(n1458) );
  CND3X2 U1740 ( .A(n3657), .B(n3658), .C(n3659), .Z(n3685) );
  CMXI2XL U1741 ( .A0(n3420), .A1(n3419), .S(n2191), .Z(n3421) );
  CMXI2XL U1742 ( .A0(n3627), .A1(n3626), .S(n2191), .Z(n3628) );
  CMXI2XL U1743 ( .A0(\reg_mem[5][16] ), .A1(\reg_mem[13][16] ), .S(net87518), 
        .Z(n3017) );
  CMXI2XL U1744 ( .A0(\reg_mem[23][16] ), .A1(\reg_mem[31][16] ), .S(net87518), 
        .Z(n3030) );
  CMXI2XL U1745 ( .A0(\reg_mem[20][17] ), .A1(\reg_mem[28][17] ), .S(net87518), 
        .Z(n2994) );
  CMXI2XL U1746 ( .A0(\reg_mem[5][14] ), .A1(\reg_mem[13][14] ), .S(net87518), 
        .Z(n3096) );
  CIVXL U1747 ( .A(net87507), .Z(n1460) );
  CMXI2XL U1748 ( .A0(\reg_mem[17][20] ), .A1(\reg_mem[25][20] ), .S(net87518), 
        .Z(n2890) );
  CNIVX2 U1749 ( .A(net87512), .Z(net87518) );
  CND2IXL U1750 ( .B(n2784), .A(n2783), .Z(N292) );
  CNR2X1 U1751 ( .A(n2664), .B(n1484), .Z(n2665) );
  CNR2X1 U1752 ( .A(n1482), .B(n1483), .Z(n1484) );
  CND2IXL U1753 ( .B(net87863), .A(n1984), .Z(n1982) );
  CND2XL U1754 ( .A(n2541), .B(n2540), .Z(n2545) );
  CND2XL U1755 ( .A(n2054), .B(n2055), .Z(n2149) );
  CMXI2XL U1756 ( .A0(n2795), .A1(n2794), .S(net87265), .Z(n2797) );
  CMXI2XL U1757 ( .A0(n3619), .A1(n3618), .S(n2199), .Z(n3620) );
  CMXI2XL U1758 ( .A0(n2933), .A1(n2932), .S(n2199), .Z(n2934) );
  CMXI2XL U1759 ( .A0(n3274), .A1(n3273), .S(n2199), .Z(n3278) );
  CMXI2XL U1760 ( .A0(\reg_mem[2][19] ), .A1(\reg_mem[10][19] ), .S(net87521), 
        .Z(n2910) );
  CNIVX1 U1761 ( .A(n1699), .Z(n1461) );
  CNIVX1 U1762 ( .A(n1463), .Z(n1462) );
  CNIVX1 U1763 ( .A(n1464), .Z(n1463) );
  CNIVX1 U1764 ( .A(regB[18]), .Z(n1464) );
  CNIVX1 U1765 ( .A(n1738), .Z(n1465) );
  CAOR2X2 U1766 ( .A(\reg_mem[9][13] ), .B(n2286), .C(n2289), .D(net83054), 
        .Z(n1074) );
  CAOR2X2 U1767 ( .A(\reg_mem[8][13] ), .B(n2280), .C(n2282), .D(n177), .Z(
        n1106) );
  CIVDX1 U1768 ( .A(prog_count_o[2]), .Z1(n1934) );
  CNIVX3 U1769 ( .A(n2078), .Z(n2096) );
  CNIVX4 U1770 ( .A(net87514), .Z(net87540) );
  CNIVX2 U1771 ( .A(net87514), .Z(net87545) );
  CNIVX4 U1772 ( .A(net87511), .Z(net87522) );
  CNIVX2 U1773 ( .A(net87374), .Z(net87391) );
  CNIVX4 U1774 ( .A(net87622), .Z(net87637) );
  CMX2XL U1775 ( .A0(n3143), .A1(n3142), .S(net87537), .Z(n1468) );
  CIVDX2 U1776 ( .A(n2169), .Z0(n1469), .Z1(n1470) );
  CND2XL U1777 ( .A(N194), .B(n3704), .Z(n2710) );
  CND2X1 U1778 ( .A(N194), .B(n2140), .Z(n2709) );
  CMXI2X1 U1779 ( .A0(n3169), .A1(n3170), .S(n2164), .Z(n3174) );
  CMXI2X1 U1780 ( .A0(\reg_mem[28][12] ), .A1(\reg_mem[24][12] ), .S(net87231), 
        .Z(n3170) );
  CND2X1 U1781 ( .A(n3003), .B(net87410), .Z(n1487) );
  CMXI2X1 U1782 ( .A0(\reg_mem[20][20] ), .A1(\reg_mem[28][20] ), .S(net87537), 
        .Z(n2887) );
  CIVXL U1783 ( .A(net87279), .Z(n1471) );
  CNIVX3 U1784 ( .A(net87235), .Z(net87247) );
  CND2IX1 U1785 ( .B(n2060), .A(net78726), .Z(n1472) );
  CND2IX1 U1786 ( .B(n2060), .A(net78726), .Z(net83575) );
  CMXI2X1 U1787 ( .A0(n4862), .A1(n4892), .S(n2096), .Z(n2679) );
  CND2XL U1788 ( .A(n1983), .B(net87863), .Z(n1985) );
  CNIVX3 U1789 ( .A(net87512), .Z(net87531) );
  CNIVX3 U1790 ( .A(net87513), .Z(net87544) );
  CNIVX3 U1791 ( .A(net87514), .Z(net87519) );
  CNIVX3 U1792 ( .A(net87514), .Z(net87529) );
  CMX2XL U1793 ( .A0(n5066), .A1(n5086), .S(n2086), .Z(n2507) );
  CMXI2X1 U1794 ( .A0(n3157), .A1(n3158), .S(n2171), .Z(n3159) );
  CMXI2X1 U1795 ( .A0(n2988), .A1(n2987), .S(net87247), .Z(n2989) );
  CND2IX1 U1796 ( .B(n1473), .A(net87230), .Z(n2130) );
  CIVX20 U1797 ( .A(\reg_mem[11][1] ), .Z(n1473) );
  CND2XL U1798 ( .A(n1985), .B(n1982), .Z(n1981) );
  CIVDX2 U1799 ( .A(net87537), .Z0(n1531), .Z1(n1532) );
  CIVX3 U1800 ( .A(n1531), .Z(net87856) );
  CMXI2XL U1801 ( .A0(n2570), .A1(n2569), .S(n2184), .Z(n2574) );
  CMXI2XL U1802 ( .A0(n2833), .A1(n2832), .S(n2184), .Z(n2834) );
  CMXI2XL U1803 ( .A0(n3045), .A1(n3044), .S(n2184), .Z(n3046) );
  CMXI2XL U1804 ( .A0(n3011), .A1(n3010), .S(n2184), .Z(n3012) );
  CMXI2XL U1805 ( .A0(n2698), .A1(n2697), .S(n2184), .Z(n2699) );
  CNIVX3 U1806 ( .A(net87235), .Z(net87248) );
  CMXI2X1 U1807 ( .A0(n2510), .A1(n2509), .S(n2197), .Z(n2511) );
  CIVX3 U1808 ( .A(n2171), .Z(n2197) );
  CMXI2X1 U1809 ( .A0(n2513), .A1(n2514), .S(n2133), .Z(n2518) );
  CMXI2X1 U1810 ( .A0(n3162), .A1(n3161), .S(n1532), .Z(n3178) );
  CND2IX2 U1811 ( .B(net87372), .A(n2158), .Z(n3671) );
  CAN2X2 U1812 ( .A(net87507), .B(net87231), .Z(n2158) );
  CIVX2 U1813 ( .A(n1474), .Z(n1476) );
  CMXI2X1 U1814 ( .A0(n2533), .A1(n2534), .S(net87508), .Z(n2535) );
  CMXI2XL U1815 ( .A0(n2999), .A1(n3000), .S(n2133), .Z(n3001) );
  CMXI2X1 U1816 ( .A0(\reg_mem[7][23] ), .A1(\reg_mem[15][23] ), .S(net87524), 
        .Z(n2756) );
  CIVX1 U1817 ( .A(n2073), .Z(n2022) );
  CIVXL U1818 ( .A(net87489), .Z(n1477) );
  CIVXL U1819 ( .A(n1477), .Z(n1478) );
  CMXI2X1 U1820 ( .A0(n3179), .A1(n3180), .S(n1482), .Z(N281) );
  CNIVX4 U1821 ( .A(net87235), .Z(net87250) );
  CMXI2XL U1822 ( .A0(n3402), .A1(n3401), .S(net87277), .Z(n3410) );
  CNR2XL U1823 ( .A(net86999), .B(n2460), .Z(n1479) );
  COND1XL U1824 ( .A(n2796), .B(n2797), .C(n3615), .Z(n2824) );
  CMXI2X1 U1825 ( .A0(\reg_mem[19][24] ), .A1(\reg_mem[3][24] ), .S(n2072), 
        .Z(n2732) );
  CNIVX4 U1826 ( .A(net87248), .Z(n1480) );
  CAN2X2 U1827 ( .A(n2163), .B(net83592), .Z(net80177) );
  CAN2XL U1828 ( .A(n1533), .B(n2711), .Z(n1481) );
  CNR2X1 U1829 ( .A(n2707), .B(n1481), .Z(n2708) );
  COND3XL U1830 ( .A(n2123), .B(n2671), .C(n2670), .D(n2669), .Z(n2711) );
  CIVXL U1831 ( .A(n1533), .Z(n1482) );
  CIVX1 U1832 ( .A(n2668), .Z(n1483) );
  CNR2IX1 U1833 ( .B(n2702), .A(n2659), .Z(n2660) );
  CND2X1 U1834 ( .A(n3004), .B(n1485), .Z(n1486) );
  CND2X1 U1835 ( .A(n1486), .B(n1487), .Z(n2064) );
  CIVXL U1836 ( .A(net87389), .Z(n1485) );
  CIVX2 U1837 ( .A(inst_fetch[1]), .Z(net78797) );
  CMXI2X1 U1838 ( .A0(n3177), .A1(n3178), .S(n2075), .Z(n3180) );
  CIVX1 U1839 ( .A(n2085), .Z(n2075) );
  CND2XL U1840 ( .A(alu_op_c[14]), .B(n1488), .Z(n1489) );
  CND2X1 U1841 ( .A(n2150), .B(n1534), .Z(n1490) );
  CND2X1 U1842 ( .A(n1490), .B(n1489), .Z(N283) );
  CIVXL U1843 ( .A(n1534), .Z(n1488) );
  CMX2X1 U1844 ( .A0(n1491), .A1(n1492), .S(n2022), .Z(n2150) );
  CMXI2XL U1845 ( .A0(n3100), .A1(n3099), .S(n2070), .Z(n1491) );
  CMXI2XL U1846 ( .A0(n3114), .A1(n3113), .S(net87389), .Z(n1492) );
  CMXI2X1 U1847 ( .A0(n3572), .A1(n3573), .S(n1496), .Z(n3580) );
  CIVX2 U1848 ( .A(net87385), .Z(n1496) );
  CMXI2X1 U1849 ( .A0(n2640), .A1(n2641), .S(n2172), .Z(n2645) );
  CMXI2X1 U1850 ( .A0(n3213), .A1(n3214), .S(n1534), .Z(N280) );
  CMXI2XL U1851 ( .A0(n3190), .A1(n3189), .S(n2176), .Z(n3194) );
  CMXI2XL U1852 ( .A0(n3542), .A1(n3541), .S(n1389), .Z(n3556) );
  CMXI2X1 U1853 ( .A0(n3102), .A1(n3101), .S(n2198), .Z(n3106) );
  CIVX3 U1854 ( .A(n2171), .Z(n2198) );
  CMXI2XL U1855 ( .A0(\reg_mem[10][27] ), .A1(\reg_mem[26][27] ), .S(n2091), 
        .Z(n2604) );
  CMXI2XL U1856 ( .A0(n5166), .A1(n5190), .S(n2091), .Z(n3678) );
  CMXI2XL U1857 ( .A0(n4667), .A1(n4697), .S(n2080), .Z(n2839) );
  CMXI2XL U1858 ( .A0(\reg_mem[8][31] ), .A1(\reg_mem[24][31] ), .S(n2080), 
        .Z(n3661) );
  CMXI2XL U1859 ( .A0(n5160), .A1(n5184), .S(n2080), .Z(n3676) );
  CMXI2XL U1860 ( .A0(\reg_mem[15][18] ), .A1(\reg_mem[31][18] ), .S(n2086), 
        .Z(n2967) );
  CMXI2X1 U1861 ( .A0(n3193), .A1(n3194), .S(n1496), .Z(n3195) );
  CMXI2X1 U1862 ( .A0(n3088), .A1(n3087), .S(n1450), .Z(n3092) );
  CIVX2 U1863 ( .A(n1493), .Z(n1495) );
  CNIVX3 U1864 ( .A(net87512), .Z(net87521) );
  CMXI2X1 U1865 ( .A0(n3195), .A1(n3196), .S(net87508), .Z(n3212) );
  CMXI2XL U1866 ( .A0(n3165), .A1(n3166), .S(n2133), .Z(n3167) );
  CMXI2X1 U1867 ( .A0(n3211), .A1(n3212), .S(n2075), .Z(n3214) );
  CND2X1 U1868 ( .A(n2990), .B(n1496), .Z(n1497) );
  CND2X1 U1869 ( .A(n2989), .B(net87385), .Z(n1498) );
  CND2X1 U1870 ( .A(n1497), .B(n1498), .Z(n2063) );
  CMXI2XL U1871 ( .A0(n2979), .A1(n2980), .S(n2172), .Z(n2981) );
  CND2IX2 U1872 ( .B(inst_fetch[3]), .A(n2013), .Z(net78798) );
  CNIVX3 U1873 ( .A(net87514), .Z(net87542) );
  CNIVX3 U1874 ( .A(n2077), .Z(n1975) );
  CNIVX3 U1875 ( .A(n2077), .Z(n2082) );
  CIVX2 U1876 ( .A(\reg_mem[10][18] ), .Z(n1542) );
  CIVX2 U1877 ( .A(\reg_mem[3][13] ), .Z(n1596) );
  CIVX2 U1878 ( .A(\reg_mem[2][13] ), .Z(n1595) );
  CIVX2 U1879 ( .A(\reg_mem[0][13] ), .Z(n1973) );
  CIVX2 U1880 ( .A(\reg_mem[10][6] ), .Z(n1965) );
  CIVX2 U1881 ( .A(\reg_mem[11][6] ), .Z(n1966) );
  CIVX2 U1882 ( .A(\reg_mem[8][6] ), .Z(n1657) );
  CIVX2 U1883 ( .A(\reg_mem[12][6] ), .Z(n1661) );
  CIVX2 U1884 ( .A(\reg_mem[10][9] ), .Z(n1601) );
  CIVX2 U1885 ( .A(\reg_mem[0][12] ), .Z(n1969) );
  CIVX2 U1886 ( .A(\reg_mem[1][12] ), .Z(n1970) );
  CIVX2 U1887 ( .A(\reg_mem[2][12] ), .Z(n1958) );
  CND2X2 U1888 ( .A(n2456), .B(n2041), .Z(n3116) );
  CNR2IX1 U1889 ( .B(N97), .A(n2270), .Z(n3558) );
  CIVX4 U1890 ( .A(n3116), .Z(n3697) );
  CIVX2 U1891 ( .A(net87243), .Z(net87230) );
  CIVX2 U1892 ( .A(inst_fetch[31]), .Z(n2043) );
  CIVX2 U1893 ( .A(inst_fetch[30]), .Z(n2060) );
  CNR2X1 U1894 ( .A(opcode_ex[1]), .B(opcode_ex[3]), .Z(n2156) );
  CIVX2 U1895 ( .A(\reg_mem[21][18] ), .Z(n1554) );
  CIVX2 U1896 ( .A(\reg_mem[20][18] ), .Z(n1553) );
  CIVX2 U1897 ( .A(\reg_mem[2][18] ), .Z(n1546) );
  CIVX2 U1898 ( .A(\reg_mem[3][18] ), .Z(n1547) );
  CIVX2 U1899 ( .A(\reg_mem[1][18] ), .Z(n1549) );
  CIVX2 U1900 ( .A(\reg_mem[0][18] ), .Z(n1548) );
  CIVX2 U1901 ( .A(\reg_mem[3][3] ), .Z(n1570) );
  CIVX2 U1902 ( .A(\reg_mem[2][3] ), .Z(n1569) );
  CIVX2 U1903 ( .A(\reg_mem[9][3] ), .Z(n1586) );
  CIVX2 U1904 ( .A(\reg_mem[8][3] ), .Z(n1585) );
  CIVX2 U1905 ( .A(\reg_mem[18][3] ), .Z(n1619) );
  CIVX2 U1906 ( .A(\reg_mem[19][3] ), .Z(n1620) );
  CIVX2 U1907 ( .A(\reg_mem[21][3] ), .Z(n1592) );
  CIVX2 U1908 ( .A(\reg_mem[20][3] ), .Z(n1591) );
  CIVX2 U1909 ( .A(\reg_mem[17][3] ), .Z(n1628) );
  CIVX2 U1910 ( .A(\reg_mem[16][3] ), .Z(n1627) );
  CIVX2 U1911 ( .A(\reg_mem[18][13] ), .Z(n1575) );
  CIVX2 U1912 ( .A(\reg_mem[19][13] ), .Z(n1576) );
  CIVX2 U1913 ( .A(\reg_mem[21][13] ), .Z(n1568) );
  CIVX2 U1914 ( .A(\reg_mem[20][13] ), .Z(n1567) );
  CIVX2 U1915 ( .A(\reg_mem[17][13] ), .Z(n1540) );
  CIVX2 U1916 ( .A(\reg_mem[16][13] ), .Z(n1539) );
  CIVX2 U1917 ( .A(\reg_mem[11][13] ), .Z(n1608) );
  CIVX2 U1918 ( .A(\reg_mem[10][13] ), .Z(n1607) );
  CIVX2 U1919 ( .A(\reg_mem[10][11] ), .Z(n1653) );
  CIVX2 U1920 ( .A(\reg_mem[11][11] ), .Z(n1654) );
  CIVX2 U1921 ( .A(\reg_mem[10][2] ), .Z(n1563) );
  CIVX2 U1922 ( .A(\reg_mem[11][2] ), .Z(n1564) );
  CIVX2 U1923 ( .A(\reg_mem[13][2] ), .Z(n2028) );
  CIVX2 U1924 ( .A(\reg_mem[12][2] ), .Z(n2027) );
  CIVX2 U1925 ( .A(\reg_mem[9][2] ), .Z(n2032) );
  CIVX2 U1926 ( .A(\reg_mem[8][2] ), .Z(n2031) );
  CIVX2 U1927 ( .A(\reg_mem[0][2] ), .Z(n1559) );
  CIVX2 U1928 ( .A(\reg_mem[1][2] ), .Z(n1560) );
  CIVX2 U1929 ( .A(\reg_mem[3][2] ), .Z(n1640) );
  CIVX2 U1930 ( .A(\reg_mem[2][2] ), .Z(n1639) );
  CIVX2 U1931 ( .A(\reg_mem[19][2] ), .Z(n1953) );
  CIVX2 U1932 ( .A(\reg_mem[18][2] ), .Z(n1952) );
  CIVX2 U1933 ( .A(\reg_mem[21][2] ), .Z(n1600) );
  CIVX2 U1934 ( .A(\reg_mem[20][2] ), .Z(n1599) );
  CIVX2 U1935 ( .A(\reg_mem[10][4] ), .Z(n1641) );
  CIVX2 U1936 ( .A(\reg_mem[11][4] ), .Z(n1642) );
  CIVX2 U1937 ( .A(\reg_mem[1][4] ), .Z(n1574) );
  CIVX2 U1938 ( .A(\reg_mem[0][4] ), .Z(n1573) );
  CIVX2 U1939 ( .A(\reg_mem[18][4] ), .Z(n1571) );
  CIVX2 U1940 ( .A(\reg_mem[19][4] ), .Z(n1572) );
  CIVX2 U1941 ( .A(\reg_mem[21][4] ), .Z(n1558) );
  CIVX2 U1942 ( .A(\reg_mem[20][4] ), .Z(n1557) );
  CIVX2 U1943 ( .A(\reg_mem[16][6] ), .Z(n1589) );
  CIVX2 U1944 ( .A(\reg_mem[17][6] ), .Z(n1590) );
  CIVX2 U1945 ( .A(\reg_mem[4][6] ), .Z(n1680) );
  CIVX2 U1946 ( .A(\reg_mem[5][6] ), .Z(n1681) );
  CIVX2 U1947 ( .A(\reg_mem[1][6] ), .Z(n1675) );
  CIVX2 U1948 ( .A(\reg_mem[0][6] ), .Z(n1674) );
  CIVX2 U1949 ( .A(\reg_mem[3][6] ), .Z(n1673) );
  CIVX2 U1950 ( .A(\reg_mem[2][6] ), .Z(n1672) );
  CIVX2 U1951 ( .A(\reg_mem[1][9] ), .Z(n1650) );
  CIVX2 U1952 ( .A(\reg_mem[0][9] ), .Z(n1649) );
  CIVX2 U1953 ( .A(\reg_mem[19][5] ), .Z(n1666) );
  CIVX2 U1954 ( .A(\reg_mem[18][5] ), .Z(n1665) );
  CIVX2 U1955 ( .A(\reg_mem[21][5] ), .Z(n1578) );
  CIVX2 U1956 ( .A(\reg_mem[20][5] ), .Z(n1577) );
  CIVX2 U1957 ( .A(\reg_mem[5][5] ), .Z(n1616) );
  CIVX2 U1958 ( .A(\reg_mem[4][5] ), .Z(n1615) );
  CIVX2 U1959 ( .A(\reg_mem[19][17] ), .Z(n1964) );
  CIVX2 U1960 ( .A(\reg_mem[18][17] ), .Z(n1963) );
  CIVX2 U1961 ( .A(\reg_mem[9][24] ), .Z(n1622) );
  CIVX2 U1962 ( .A(\reg_mem[8][24] ), .Z(n1621) );
  CIVX2 U1963 ( .A(\reg_mem[13][24] ), .Z(n1562) );
  CIVX2 U1964 ( .A(\reg_mem[12][24] ), .Z(n1561) );
  CIVX2 U1965 ( .A(\reg_mem[2][24] ), .Z(n1587) );
  CIVX2 U1966 ( .A(\reg_mem[3][24] ), .Z(n1588) );
  CIVX2 U1967 ( .A(\reg_mem[5][24] ), .Z(n1584) );
  CIVX2 U1968 ( .A(\reg_mem[4][24] ), .Z(n1583) );
  CIVX2 U1969 ( .A(\reg_mem[1][24] ), .Z(n1626) );
  CIVX2 U1970 ( .A(\reg_mem[0][24] ), .Z(n1625) );
  CIVX2 U1971 ( .A(\reg_mem[17][24] ), .Z(n1671) );
  CIVX2 U1972 ( .A(\reg_mem[16][24] ), .Z(n1670) );
  CIVX2 U1973 ( .A(\reg_mem[19][24] ), .Z(n1636) );
  CIVX2 U1974 ( .A(\reg_mem[18][24] ), .Z(n1635) );
  CIVX2 U1975 ( .A(\reg_mem[21][24] ), .Z(n1955) );
  CIVX2 U1976 ( .A(\reg_mem[20][24] ), .Z(n1954) );
  CIVX2 U1977 ( .A(\reg_mem[9][28] ), .Z(n1679) );
  CIVX2 U1978 ( .A(\reg_mem[8][28] ), .Z(n1678) );
  CIVX2 U1979 ( .A(\reg_mem[13][28] ), .Z(n1949) );
  CIVX2 U1980 ( .A(\reg_mem[12][28] ), .Z(n1948) );
  CIVX2 U1981 ( .A(\reg_mem[9][31] ), .Z(n1566) );
  CIVX2 U1982 ( .A(\reg_mem[8][31] ), .Z(n1565) );
  CIVX2 U1983 ( .A(\reg_mem[13][31] ), .Z(n1582) );
  CIVX2 U1984 ( .A(\reg_mem[12][31] ), .Z(n1581) );
  CIVX2 U1985 ( .A(\reg_mem[0][27] ), .Z(n1971) );
  CIVX2 U1986 ( .A(\reg_mem[1][27] ), .Z(n1972) );
  CIVX2 U1987 ( .A(\reg_mem[9][27] ), .Z(n1614) );
  CIVX2 U1988 ( .A(\reg_mem[8][27] ), .Z(n1613) );
  CIVX2 U1989 ( .A(\reg_mem[11][27] ), .Z(n1606) );
  CIVX2 U1990 ( .A(\reg_mem[10][27] ), .Z(n1605) );
  CIVX2 U1991 ( .A(\reg_mem[13][27] ), .Z(n1656) );
  CIVX2 U1992 ( .A(\reg_mem[12][27] ), .Z(n1655) );
  CIVX2 U1993 ( .A(\reg_mem[19][27] ), .Z(n1664) );
  CIVX2 U1994 ( .A(\reg_mem[18][27] ), .Z(n1663) );
  CIVX2 U1995 ( .A(\reg_mem[16][27] ), .Z(n1629) );
  CIVX2 U1996 ( .A(\reg_mem[17][27] ), .Z(n1630) );
  CIVX2 U1997 ( .A(\reg_mem[21][27] ), .Z(n1550) );
  CIVX2 U1998 ( .A(\reg_mem[20][27] ), .Z(n1551) );
  CIVX2 U1999 ( .A(\reg_mem[5][19] ), .Z(n1648) );
  CIVX2 U2000 ( .A(\reg_mem[4][19] ), .Z(n1647) );
  CIVX2 U2001 ( .A(\reg_mem[21][19] ), .Z(n1598) );
  CIVX2 U2002 ( .A(\reg_mem[20][19] ), .Z(n1597) );
  CIVX2 U2003 ( .A(\reg_mem[8][20] ), .Z(n1611) );
  CIVX2 U2004 ( .A(\reg_mem[9][20] ), .Z(n1612) );
  CIVX2 U2005 ( .A(\reg_mem[5][0] ), .Z(n1593) );
  CIVX2 U2006 ( .A(\reg_mem[17][0] ), .Z(n1644) );
  CIVX2 U2007 ( .A(\reg_mem[16][0] ), .Z(n1643) );
  CIVX2 U2008 ( .A(\reg_mem[21][0] ), .Z(n1660) );
  CIVX2 U2009 ( .A(\reg_mem[20][0] ), .Z(n1659) );
  CIVX2 U2010 ( .A(\reg_mem[10][0] ), .Z(n1617) );
  CIVX2 U2011 ( .A(\reg_mem[11][0] ), .Z(n1618) );
  CIVX2 U2012 ( .A(\reg_mem[2][7] ), .Z(n1609) );
  CIVX2 U2013 ( .A(\reg_mem[3][7] ), .Z(n1610) );
  CIVX2 U2014 ( .A(\reg_mem[9][7] ), .Z(n1646) );
  CIVX2 U2015 ( .A(\reg_mem[8][7] ), .Z(n1645) );
  CIVX2 U2016 ( .A(\reg_mem[17][7] ), .Z(n1638) );
  CIVX2 U2017 ( .A(\reg_mem[16][7] ), .Z(n1637) );
  CIVX2 U2018 ( .A(\reg_mem[18][10] ), .Z(n1544) );
  CIVX2 U2019 ( .A(\reg_mem[19][10] ), .Z(n1545) );
  CIVX2 U2020 ( .A(\reg_mem[8][8] ), .Z(n1633) );
  CIVX2 U2021 ( .A(\reg_mem[9][8] ), .Z(n1634) );
  CIVX2 U2022 ( .A(\reg_mem[11][8] ), .Z(n1962) );
  CIVX2 U2023 ( .A(\reg_mem[10][8] ), .Z(n1961) );
  CIVX2 U2024 ( .A(\reg_mem[2][8] ), .Z(n1631) );
  CIVX2 U2025 ( .A(\reg_mem[3][8] ), .Z(n1632) );
  CIVX2 U2026 ( .A(\reg_mem[19][8] ), .Z(n1652) );
  CIVX2 U2027 ( .A(\reg_mem[18][8] ), .Z(n1651) );
  CIVX2 U2028 ( .A(\reg_mem[4][12] ), .Z(n1676) );
  CIVX2 U2029 ( .A(\reg_mem[5][12] ), .Z(n1677) );
  CIVX2 U2030 ( .A(\reg_mem[20][12] ), .Z(n1579) );
  CIVX2 U2031 ( .A(\reg_mem[21][12] ), .Z(n1580) );
  CIVX2 U2032 ( .A(\reg_mem[9][12] ), .Z(n1951) );
  CIVX2 U2033 ( .A(\reg_mem[8][12] ), .Z(n1950) );
  CIVX2 U2034 ( .A(\reg_mem[11][12] ), .Z(n1624) );
  CIVX2 U2035 ( .A(\reg_mem[10][12] ), .Z(n1623) );
  CIVX2 U2036 ( .A(\reg_mem[13][12] ), .Z(n1604) );
  CIVX2 U2037 ( .A(\reg_mem[12][12] ), .Z(n1603) );
  CNR2XL U2038 ( .A(n2115), .B(n2620), .Z(n2621) );
  CNR2IXL U2039 ( .B(N122), .A(n2271), .Z(n2630) );
  CNR3X1 U2040 ( .A(n5267), .B(n230), .C(n5266), .Z(n198) );
  CND3XL U2041 ( .A(n194), .B(n1939), .C(n210), .Z(n211) );
  CNR2IX1 U2042 ( .B(n207), .A(n208), .Z(n219) );
  CNIVX2 U2043 ( .A(data_mem_rd_d), .Z(n2202) );
  CIVX2 U2044 ( .A(\reg_mem[11][18] ), .Z(n1543) );
  CIVX2 U2045 ( .A(\reg_mem[1][13] ), .Z(n1974) );
  CIVX2 U2046 ( .A(\reg_mem[9][6] ), .Z(n1658) );
  CIVX2 U2047 ( .A(\reg_mem[13][6] ), .Z(n1662) );
  CIVX2 U2048 ( .A(\reg_mem[11][9] ), .Z(n1602) );
  CIVX2 U2049 ( .A(net86657), .Z(net87990) );
  CIVX2 U2050 ( .A(\reg_mem[3][12] ), .Z(n1959) );
  CNR3XL U2051 ( .A(n3076), .B(n3075), .C(n3074), .Z(n3077) );
  CNR3XL U2052 ( .A(n2862), .B(n2863), .C(n2864), .Z(n2865) );
  CND3XL U2053 ( .A(n2855), .B(n2854), .C(n2853), .Z(n2863) );
  CNR2IXL U2054 ( .B(N112), .A(n2115), .Z(n3005) );
  CNR2IXL U2055 ( .B(N108), .A(n2271), .Z(n3146) );
  CNR2IXL U2056 ( .B(N105), .A(n2123), .Z(n3250) );
  CND2X1 U2057 ( .A(n3637), .B(n3636), .Z(n3643) );
  CND2X1 U2058 ( .A(n3524), .B(n3523), .Z(alu_op_c[2]) );
  CANR1X1 U2059 ( .A(N65), .B(n3697), .C(n3560), .Z(n3561) );
  CNR2IX1 U2060 ( .B(n3559), .A(n3558), .Z(n3562) );
  CIVDX1 U2061 ( .A(n201), .Z0(n1500), .Z1(n1501) );
  CIVX2 U2062 ( .A(n193), .Z(n2431) );
  CIVDX1 U2063 ( .A(n199), .Z0(n1502), .Z1(n1503) );
  CND2X1 U2064 ( .A(n228), .B(n194), .Z(n232) );
  COND3X1 U2065 ( .A(data_mem_rd_d), .B(n2213), .C(n206), .D(n228), .Z(n238)
         );
  CIVDX1 U2066 ( .A(n216), .Z0(n1504), .Z1(n1505) );
  CIVDX1 U2067 ( .A(n215), .Z0(n1506), .Z1(n1507) );
  CND3X1 U2068 ( .A(n191), .B(n1939), .C(n202), .Z(n201) );
  CIVDX1 U2069 ( .A(n217), .Z0(n1508), .Z1(n1509) );
  CIVDX1 U2070 ( .A(n205), .Z0(n1510), .Z1(n1511) );
  CIVDX1 U2071 ( .A(n203), .Z0(n1512), .Z1(n1513) );
  CIVDX1 U2072 ( .A(n197), .Z0(n1514), .Z1(n1515) );
  CND3X1 U2073 ( .A(n206), .B(n1939), .C(n210), .Z(n217) );
  CND3X1 U2074 ( .A(n204), .B(n1939), .C(n210), .Z(n216) );
  CND3X1 U2075 ( .A(n202), .B(n1939), .C(n210), .Z(n215) );
  CND3XL U2076 ( .A(n198), .B(n1939), .C(n219), .Z(n222) );
  CND3XL U2077 ( .A(n196), .B(n1939), .C(n219), .Z(n221) );
  CND3XL U2078 ( .A(n192), .B(n1939), .C(n219), .Z(n218) );
  CND3X1 U2079 ( .A(n200), .B(n1939), .C(n219), .Z(n223) );
  CND2XL U2080 ( .A(n196), .B(n191), .Z(n195) );
  CND2XL U2081 ( .A(n194), .B(n191), .Z(n193) );
  CND2XL U2082 ( .A(n191), .B(n192), .Z(n158) );
  CIVDX1 U2083 ( .A(n214), .Z0(n1516), .Z1(n1517) );
  CND3X1 U2084 ( .A(n200), .B(n1939), .C(n210), .Z(n214) );
  CIVDX1 U2085 ( .A(n213), .Z0(n1518), .Z1(n1519) );
  CND3X1 U2086 ( .A(n198), .B(n1939), .C(n210), .Z(n213) );
  CIVDX1 U2087 ( .A(n212), .Z0(n1520), .Z1(n1521) );
  CND3X1 U2088 ( .A(n196), .B(n1939), .C(n210), .Z(n212) );
  CND3X1 U2089 ( .A(n191), .B(n1939), .C(n206), .Z(n205) );
  CND3X1 U2090 ( .A(n191), .B(n1939), .C(n204), .Z(n203) );
  CIVX2 U2091 ( .A(n199), .Z(n2404) );
  CIVX2 U2092 ( .A(n197), .Z(n2410) );
  CIVDX1 U2093 ( .A(n224), .Z0(n1522), .Z1(n1523) );
  CND3X1 U2094 ( .A(n191), .B(n1939), .C(n200), .Z(n199) );
  CND3X1 U2095 ( .A(n191), .B(n1939), .C(n198), .Z(n197) );
  CND2XL U2096 ( .A(n228), .B(n196), .Z(n233) );
  CIVDX1 U2097 ( .A(n224), .Z0(n1524), .Z1(n1525) );
  CIVDX1 U2098 ( .A(n220), .Z0(n1526), .Z1(n1527) );
  CND3X1 U2099 ( .A(n194), .B(n1939), .C(n219), .Z(n220) );
  CIVDX1 U2100 ( .A(n211), .Z0(n1528), .Z1(n1529) );
  CIVDX1 U2101 ( .A(n238), .Z1(n1530) );
  CND2XL U2102 ( .A(n228), .B(n202), .Z(n236) );
  CND3X1 U2103 ( .A(n202), .B(n1939), .C(n219), .Z(n224) );
  CND2XL U2104 ( .A(n228), .B(n198), .Z(n234) );
  CIVX2 U2105 ( .A(net79756), .Z(net87374) );
  CNIVX2 U2106 ( .A(net87379), .Z(net87408) );
  CIVX2 U2107 ( .A(net87400), .Z(net87483) );
  CIVX2 U2108 ( .A(n2167), .Z(n2169) );
  CIVX2 U2109 ( .A(net87799), .Z(n1993) );
  CIVDX4 U2110 ( .A(n3615), .Z0(n1533), .Z1(n1534) );
  CIVXL U2111 ( .A(opcode_ex[3]), .Z(n2450) );
  CAN2X1 U2112 ( .A(n2121), .B(n2122), .Z(n1536) );
  CAN2X1 U2113 ( .A(n2130), .B(n2131), .Z(n1537) );
  CAOR2X1 U2114 ( .A(N140), .B(n3701), .C(n3476), .D(n3475), .Z(n1538) );
  CND4XL U2115 ( .A(i_type), .B(immi_val[31]), .C(n5239), .D(n2441), .Z(n3286)
         );
  CIVX4 U2116 ( .A(n2164), .Z(n2165) );
  CIVX2 U2117 ( .A(n2172), .Z(n2185) );
  CMXI2XL U2118 ( .A0(n1539), .A1(n1540), .S(net87797), .Z(n4304) );
  CIVX1 U2119 ( .A(alu_op_c[19]), .Z(n2940) );
  CMXI2XL U2120 ( .A0(n4995), .A1(n4996), .S(net88175), .Z(n5022) );
  CMXI2X1 U2121 ( .A0(n4099), .A1(n4100), .S(n1988), .Z(n4101) );
  CIVX1 U2122 ( .A(n3563), .Z(n3741) );
  CIVXL U2123 ( .A(immi_val[0]), .Z(n1541) );
  CMXI2XL U2124 ( .A0(n3896), .A1(n3895), .S(net87628), .Z(n3902) );
  CMXI2XL U2125 ( .A0(n4096), .A1(n4095), .S(net87628), .Z(n4102) );
  CMXI2XL U2126 ( .A0(n1542), .A1(n1543), .S(net87794), .Z(n4527) );
  CMXI2XL U2127 ( .A0(n1544), .A1(n1545), .S(net87795), .Z(n4193) );
  CANR2X1 U2128 ( .A(regc_addr_wb[2]), .B(n240), .C(regb_addr_wb[2]), .D(n2116), .Z(n230) );
  CMXI2XL U2129 ( .A0(n2634), .A1(n2633), .S(n2188), .Z(n2638) );
  CND3X1 U2130 ( .A(n3290), .B(n3289), .C(n3288), .Z(alu_op_c[7]) );
  CND2IXL U2131 ( .B(n2587), .A(n2586), .Z(alu_op_c[28]) );
  CIVX2 U2132 ( .A(n2167), .Z(n2168) );
  CND2IXL U2133 ( .B(n2668), .A(n2667), .Z(alu_op_c[26]) );
  CND2XL U2134 ( .A(N195), .B(n3704), .Z(n2667) );
  CND2XL U2135 ( .A(net87642), .B(n1989), .Z(n1986) );
  CMXI2XL U2136 ( .A0(n4962), .A1(n4961), .S(net87636), .Z(n4963) );
  CMXI2XL U2137 ( .A0(n4744), .A1(n4743), .S(net87636), .Z(n4752) );
  CMXI2XL U2138 ( .A0(n4322), .A1(n4321), .S(net87635), .Z(n4323) );
  CMXI2XL U2139 ( .A0(n4520), .A1(n4519), .S(net87635), .Z(n4526) );
  CMXI2XL U2140 ( .A0(n4852), .A1(n4851), .S(net87642), .Z(n4853) );
  CMXI2XL U2141 ( .A0(n4088), .A1(n4087), .S(net87642), .Z(n4094) );
  CMXI2XL U2142 ( .A0(n4846), .A1(n4845), .S(net87642), .Z(n4854) );
  CMXI2X1 U2143 ( .A0(n2922), .A1(n2923), .S(net87483), .Z(n2939) );
  CND2X1 U2144 ( .A(net87372), .B(n2158), .Z(n3681) );
  CMXI2XL U2145 ( .A0(n1546), .A1(n1547), .S(net87806), .Z(n4519) );
  CMXI2XL U2146 ( .A0(n1548), .A1(n1549), .S(net87807), .Z(n4520) );
  CMXI2XL U2147 ( .A0(n1551), .A1(n1550), .S(net87798), .Z(n5002) );
  CND3X1 U2148 ( .A(i_type), .B(n3344), .C(n2455), .Z(n1552) );
  CND3XL U2149 ( .A(i_type), .B(n3344), .C(n2455), .Z(n3695) );
  CND2IX1 U2150 ( .B(net87404), .A(n2148), .Z(n3663) );
  CMXI2XL U2151 ( .A0(n1553), .A1(n1554), .S(net87794), .Z(n4542) );
  CMXI2X1 U2152 ( .A0(n4559), .A1(n4560), .S(n1960), .Z(n4561) );
  CMXI2XL U2153 ( .A0(n2000), .A1(net77974), .S(net87637), .Z(net77965) );
  CMXI2XL U2154 ( .A0(n4816), .A1(n4815), .S(net87637), .Z(n4822) );
  CMXI2XL U2155 ( .A0(n4824), .A1(n4823), .S(net87637), .Z(n4830) );
  CMXI2XL U2156 ( .A0(n4406), .A1(n4405), .S(net87637), .Z(n4414) );
  COND1X1 U2157 ( .A(n2154), .B(n3563), .C(enable), .Z(n2138) );
  CMXI2XL U2158 ( .A0(n3408), .A1(n3407), .S(net87256), .Z(n3409) );
  CMXI2XL U2159 ( .A0(n3404), .A1(n3403), .S(n2166), .Z(n3408) );
  CNIVX2 U2160 ( .A(net87380), .Z(net87409) );
  CNIVX2 U2161 ( .A(net87380), .Z(net87410) );
  CMXI2XL U2162 ( .A0(n3968), .A1(n3967), .S(net87725), .Z(n3969) );
  CMXI2XL U2163 ( .A0(n3970), .A1(n3969), .S(net82859), .Z(n3996) );
  CAN2XL U2164 ( .A(N191), .B(n2140), .Z(n2144) );
  CAN2X2 U2165 ( .A(n3704), .B(n1533), .Z(n2140) );
  CANR2XL U2166 ( .A(N192), .B(n2140), .C(n1533), .D(n2786), .Z(n2783) );
  CANR2XL U2167 ( .A(N189), .B(n2140), .C(n1533), .D(n2906), .Z(n2903) );
  CND2XL U2168 ( .A(N196), .B(n2140), .Z(n2624) );
  CIVXL U2169 ( .A(n2273), .Z(n2270) );
  CIVX2 U2170 ( .A(n2273), .Z(n2272) );
  CMXI2XL U2171 ( .A0(n3377), .A1(n3378), .S(n2075), .Z(n3380) );
  CIVX1 U2172 ( .A(net87405), .Z(net87372) );
  CIVX1 U2173 ( .A(net87391), .Z(net87368) );
  CMXI2XL U2174 ( .A0(n3563), .A1(enable), .S(prog_count_o[2]), .Z(n3525) );
  CIVXL U2175 ( .A(immi_val[7]), .Z(n1555) );
  CIVX2 U2176 ( .A(net78790), .Z(net87787) );
  CIVX2 U2177 ( .A(net78790), .Z(net87789) );
  CIVX2 U2178 ( .A(net78790), .Z(net87788) );
  CIVX2 U2179 ( .A(net78790), .Z(net87786) );
  CMXI2X1 U2180 ( .A0(n4535), .A1(n4536), .S(n1960), .Z(n4562) );
  CMXI2XL U2181 ( .A0(alu_op_c[2]), .A1(n3555), .S(n3615), .Z(n3557) );
  CNIVX12 U2182 ( .A(net87788), .Z(net87790) );
  CIVXL U2183 ( .A(n3481), .Z(n3482) );
  CIVXL U2184 ( .A(alu_op_c[16]), .Z(n3038) );
  CMXI2XL U2185 ( .A0(n4252), .A1(n4251), .S(net87638), .Z(n4258) );
  CMXI2XL U2186 ( .A0(n4288), .A1(n4287), .S(net87638), .Z(n4289) );
  CMXI2XL U2187 ( .A0(n3966), .A1(n3965), .S(net87638), .Z(n3967) );
  CMXI2XL U2188 ( .A0(n4688), .A1(n4687), .S(net87638), .Z(n4689) );
  CNIVX2 U2189 ( .A(net87374), .Z(net87388) );
  CNIVX2 U2190 ( .A(net87374), .Z(net87386) );
  CMXI2XL U2191 ( .A0(n4162), .A1(n4161), .S(net87627), .Z(n4170) );
  CMXI2XL U2192 ( .A0(n4078), .A1(n4077), .S(net87627), .Z(n4079) );
  CMXI2XL U2193 ( .A0(n5202), .A1(n5201), .S(net87627), .Z(n5210) );
  CMXI2XL U2194 ( .A0(n3780), .A1(n3779), .S(net87627), .Z(n3781) );
  CMXI2XL U2195 ( .A0(n4282), .A1(n4281), .S(net87627), .Z(n4290) );
  CIVXL U2196 ( .A(immi_val[5]), .Z(n1556) );
  CMXI2XL U2197 ( .A0(\reg_mem[2][3] ), .A1(\reg_mem[3][3] ), .S(n2068), .Z(
        n3488) );
  CMXI2XL U2198 ( .A0(\reg_mem[12][0] ), .A1(\reg_mem[13][0] ), .S(n2069), .Z(
        n2471) );
  CMXI2XL U2199 ( .A0(\reg_mem[18][11] ), .A1(\reg_mem[19][11] ), .S(n1456), 
        .Z(n3197) );
  CMXI2XL U2200 ( .A0(\reg_mem[4][7] ), .A1(\reg_mem[5][7] ), .S(n2070), .Z(
        n3294) );
  CMXI2XL U2201 ( .A0(\reg_mem[8][9] ), .A1(\reg_mem[9][9] ), .S(n2069), .Z(
        n3260) );
  CMXI2XL U2202 ( .A0(n3501), .A1(n3500), .S(n1532), .Z(n3517) );
  CMXI2XL U2203 ( .A0(n3493), .A1(n3492), .S(net87273), .Z(n3501) );
  CND2XL U2204 ( .A(N190), .B(n3704), .Z(n2868) );
  CMXI2XL U2205 ( .A0(n4655), .A1(n4685), .S(n2087), .Z(n2832) );
  CNR2XL U2206 ( .A(n2865), .B(n2127), .Z(n2866) );
  CMXI2XL U2207 ( .A0(n3422), .A1(n3421), .S(net87278), .Z(n3423) );
  CMXI2XL U2208 ( .A0(n3424), .A1(n3423), .S(n1389), .Z(n3425) );
  CMXI2X1 U2209 ( .A0(n2684), .A1(n2683), .S(net87280), .Z(n2685) );
  CMXI2XL U2210 ( .A0(n3135), .A1(n3134), .S(net87398), .Z(n3143) );
  CND2IX2 U2211 ( .B(n2001), .A(net87488), .Z(net78790) );
  CMXI2XL U2212 ( .A0(n1557), .A1(n1558), .S(net87797), .Z(net78495) );
  CMXI2XL U2213 ( .A0(n1559), .A1(n1560), .S(net87790), .Z(n3846) );
  CMXI2X1 U2214 ( .A0(n5001), .A1(n5002), .S(n1988), .Z(n5003) );
  CMXI2XL U2215 ( .A0(n4860), .A1(n4890), .S(n2080), .Z(n2680) );
  CMXI2X1 U2216 ( .A0(n2642), .A1(n2643), .S(n2039), .Z(n2644) );
  CMXI2X1 U2217 ( .A0(net78496), .A1(net78495), .S(n1988), .Z(net78494) );
  CMXI2XL U2218 ( .A0(n1561), .A1(n1562), .S(net87794), .Z(n4828) );
  CMXI2XL U2219 ( .A0(n1563), .A1(n1564), .S(net87790), .Z(n3853) );
  CMXI2XL U2220 ( .A0(n1565), .A1(n1566), .S(net87804), .Z(n5174) );
  CMXI2XL U2221 ( .A0(n1567), .A1(n1568), .S(net87802), .Z(n4308) );
  CMXI2XL U2222 ( .A0(n1569), .A1(n1570), .S(net87793), .Z(n3877) );
  CMXI2XL U2223 ( .A0(n1571), .A1(n1572), .S(net87790), .Z(net78502) );
  CMXI2X1 U2224 ( .A0(n4827), .A1(n4828), .S(n1988), .Z(n4829) );
  CMXI2X1 U2225 ( .A0(n5173), .A1(n5174), .S(n1988), .Z(n5180) );
  CMXI2XL U2226 ( .A0(n1573), .A1(n1574), .S(net87806), .Z(n3922) );
  CNR2IX2 U2227 ( .B(n2702), .A(n2701), .Z(n2703) );
  CMXI2XL U2228 ( .A0(n1575), .A1(n1576), .S(net87799), .Z(n4303) );
  CMXI2XL U2229 ( .A0(n1577), .A1(n1578), .S(net87803), .Z(n3976) );
  CMXI2X1 U2230 ( .A0(n3921), .A1(n3922), .S(n1988), .Z(n3928) );
  CMXI2X1 U2231 ( .A0(n4325), .A1(n4326), .S(net88175), .Z(net77918) );
  CMXI2X1 U2232 ( .A0(n3975), .A1(n3976), .S(n1988), .Z(n3977) );
  CNIVX3 U2233 ( .A(net87618), .Z(net87623) );
  CIVX12 U2234 ( .A(net87637), .Z(n1988) );
  CMXI2X1 U2235 ( .A0(\reg_mem[2][8] ), .A1(\reg_mem[3][8] ), .S(net87394), 
        .Z(n3708) );
  CMXI2X1 U2236 ( .A0(n1579), .A1(n1580), .S(net87799), .Z(n4274) );
  CMXI2XL U2237 ( .A0(n1581), .A1(n1582), .S(net87800), .Z(n5178) );
  CNR2X1 U2238 ( .A(n2115), .B(n3634), .Z(n3635) );
  CMXI2X1 U2239 ( .A0(n3283), .A1(n3284), .S(n3615), .Z(N278) );
  CMXI2XL U2240 ( .A0(n1583), .A1(n1584), .S(net87809), .Z(n4820) );
  CMXI2XL U2241 ( .A0(n1585), .A1(n1586), .S(net87794), .Z(n3886) );
  CND2X1 U2242 ( .A(n3704), .B(N200), .Z(n2137) );
  CMXI2XL U2243 ( .A0(n1587), .A1(n1588), .S(net87807), .Z(n4815) );
  CMXI2XL U2244 ( .A0(n1589), .A1(n1590), .S(net87798), .Z(n4016) );
  CMXI2XL U2245 ( .A0(n1591), .A1(n1592), .S(net87791), .Z(n3900) );
  CIVX2 U2246 ( .A(n2068), .Z(n2066) );
  CAN2XL U2247 ( .A(n1533), .B(n2869), .Z(n2127) );
  CND2IXL U2248 ( .B(n2869), .A(n2868), .Z(n5244) );
  CND2X1 U2249 ( .A(n2831), .B(n2830), .Z(n2869) );
  CMXI2XL U2250 ( .A0(n1594), .A1(n1593), .S(net87794), .Z(n3762) );
  CMXI2X1 U2251 ( .A0(n4063), .A1(n4064), .S(n1988), .Z(n4065) );
  CMXI2XL U2252 ( .A0(n1595), .A1(n1596), .S(net87795), .Z(net77974) );
  CMXI2XL U2253 ( .A0(n1597), .A1(n1598), .S(net87790), .Z(n4582) );
  CMXI2XL U2254 ( .A0(n1599), .A1(n1600), .S(net87790), .Z(net78619) );
  CND2IXL U2255 ( .B(n3081), .A(n3080), .Z(n5243) );
  CIVXL U2256 ( .A(n3612), .Z(n2686) );
  CMXI2XL U2257 ( .A0(n1601), .A1(n1602), .S(net87806), .Z(n4139) );
  CMXI2XL U2258 ( .A0(n1603), .A1(n1604), .S(net87802), .Z(n4264) );
  CMXI2XL U2259 ( .A0(n1605), .A1(n1606), .S(net87790), .Z(n4987) );
  CMXI2X1 U2260 ( .A0(n4091), .A1(n4092), .S(n1988), .Z(n4093) );
  CMXI2XL U2261 ( .A0(n1607), .A1(n1608), .S(net87795), .Z(n4295) );
  CMXI2XL U2262 ( .A0(n1609), .A1(n1610), .S(net87798), .Z(n4041) );
  CMXI2XL U2263 ( .A0(n2801), .A1(n2800), .S(n2180), .Z(n2802) );
  CMXI2XL U2264 ( .A0(n2605), .A1(n2604), .S(n2194), .Z(n2609) );
  CMXI2XL U2265 ( .A0(n2845), .A1(n2844), .S(n2194), .Z(n2846) );
  CMXI2XL U2266 ( .A0(n3661), .A1(n3660), .S(n2194), .Z(n3662) );
  CMXI2XL U2267 ( .A0(n3023), .A1(n3022), .S(n2194), .Z(n3027) );
  CMXI2X1 U2268 ( .A0(n4615), .A1(n4616), .S(n1988), .Z(n4617) );
  CMXI2XL U2269 ( .A0(n1611), .A1(n1612), .S(net87799), .Z(n4612) );
  CMXI2X1 U2270 ( .A0(n4581), .A1(n4582), .S(net88166), .Z(n4583) );
  CIVX1 U2271 ( .A(n2113), .Z(n2745) );
  CMXI2X1 U2272 ( .A0(n4015), .A1(n4016), .S(n1988), .Z(n4022) );
  CMXI2XL U2273 ( .A0(n1613), .A1(n1614), .S(net87803), .Z(n4988) );
  CMXI2X1 U2274 ( .A0(n3239), .A1(n3238), .S(n2198), .Z(n3243) );
  CIVXL U2275 ( .A(alu_op_c[10]), .Z(n3248) );
  CMXI2XL U2276 ( .A0(n1615), .A1(n1616), .S(net87795), .Z(n3958) );
  CMXI2XL U2277 ( .A0(n3575), .A1(n3574), .S(n2201), .Z(n3578) );
  CMXI2X1 U2278 ( .A0(n4599), .A1(n4600), .S(n1960), .Z(n4601) );
  CMXI2X1 U2279 ( .A0(n4987), .A1(n4988), .S(n1988), .Z(n4994) );
  CMXI2XL U2280 ( .A0(n1617), .A1(n1618), .S(net87800), .Z(n3765) );
  CMXI2XL U2281 ( .A0(n1619), .A1(n1620), .S(net87793), .Z(n3895) );
  CMXI2XL U2282 ( .A0(\reg_mem[21][14] ), .A1(\reg_mem[29][14] ), .S(net87537), 
        .Z(n3110) );
  CMXI2XL U2283 ( .A0(n1621), .A1(n1622), .S(net87791), .Z(n4824) );
  CMXI2XL U2284 ( .A0(n1623), .A1(n1624), .S(net87804), .Z(n4259) );
  CMXI2XL U2285 ( .A0(n1625), .A1(n1626), .S(net87809), .Z(n4816) );
  CMXI2XL U2286 ( .A0(n1627), .A1(n1628), .S(net87807), .Z(n3896) );
  CMXI2XL U2287 ( .A0(n1629), .A1(n1630), .S(net87798), .Z(n4998) );
  CMXI2XL U2288 ( .A0(n3426), .A1(n3425), .S(n2091), .Z(n3428) );
  CMXI2XL U2289 ( .A0(n4379), .A1(n4409), .S(n2088), .Z(n3044) );
  CMXI2XL U2290 ( .A0(n1631), .A1(n1632), .S(net87790), .Z(n4087) );
  CMXI2XL U2291 ( .A0(n1633), .A1(n1634), .S(net87799), .Z(n4096) );
  CMXI2XL U2292 ( .A0(n1635), .A1(n1636), .S(net87790), .Z(n4833) );
  CMXI2XL U2293 ( .A0(n1637), .A1(n1638), .S(net87790), .Z(n4060) );
  CMXI2X1 U2294 ( .A0(n2682), .A1(n2681), .S(n2187), .Z(n2683) );
  CMXI2XL U2295 ( .A0(n1639), .A1(n1640), .S(net87795), .Z(n3845) );
  CMXI2XL U2296 ( .A0(n1641), .A1(n1642), .S(net87795), .Z(n3929) );
  CMXI2XL U2297 ( .A0(n3109), .A1(n3110), .S(n2038), .Z(n3111) );
  CMXI2X1 U2298 ( .A0(n4609), .A1(n4610), .S(net87698), .Z(n4620) );
  CMXI2X1 U2299 ( .A0(n4301), .A1(n4302), .S(net87701), .Z(net77950) );
  CMXI2X1 U2300 ( .A0(n3321), .A1(n3322), .S(n3615), .Z(N276) );
  CMXI2XL U2301 ( .A0(n1643), .A1(n1644), .S(net87793), .Z(n3776) );
  CMXI2XL U2302 ( .A0(n1645), .A1(n1646), .S(net87791), .Z(n4050) );
  CMXI2XL U2303 ( .A0(n1647), .A1(n1648), .S(net87803), .Z(n4568) );
  CANR1X1 U2304 ( .A(N71), .B(n3697), .C(n3287), .Z(n3288) );
  CMXI2XL U2305 ( .A0(n1649), .A1(n1650), .S(net87794), .Z(n4132) );
  CMXI2XL U2306 ( .A0(n1651), .A1(n1652), .S(net87800), .Z(n4105) );
  CMXI2XL U2307 ( .A0(n1653), .A1(n1654), .S(net87806), .Z(n4219) );
  CMXI2X1 U2308 ( .A0(n4567), .A1(n4568), .S(n1988), .Z(n4569) );
  CMXI2XL U2309 ( .A0(n1655), .A1(n1656), .S(net87799), .Z(n4992) );
  CMXI2X1 U2310 ( .A0(n4131), .A1(n4132), .S(n1988), .Z(n4138) );
  CMXI2XL U2311 ( .A0(n1657), .A1(n1658), .S(net87802), .Z(n4006) );
  CMXI2XL U2312 ( .A0(n1659), .A1(n1660), .S(net87804), .Z(n3780) );
  CMXI2X1 U2313 ( .A0(n4627), .A1(n4628), .S(net87701), .Z(n4644) );
  CMXI2X1 U2314 ( .A0(n4643), .A1(n4644), .S(n1960), .Z(n4645) );
  CMXI2X1 U2315 ( .A0(net78073), .A1(net78074), .S(net82863), .Z(net78041) );
  CMXI2XL U2316 ( .A0(n1661), .A1(n1662), .S(net87798), .Z(n4010) );
  CMXI2X1 U2317 ( .A0(n4991), .A1(n4992), .S(n1988), .Z(n4993) );
  CMXI2X1 U2318 ( .A0(n4005), .A1(n4006), .S(n1988), .Z(n4012) );
  CMXI2X1 U2319 ( .A0(n4569), .A1(n4570), .S(net87699), .Z(n4578) );
  CNR2IX1 U2320 ( .B(n2134), .A(n1669), .Z(n1668) );
  CMXI2XL U2321 ( .A0(n5158), .A1(n5157), .S(net86657), .Z(N202) );
  CMXI2XL U2322 ( .A0(n4342), .A1(n4341), .S(net87717), .Z(n4343) );
  CMXI2X1 U2323 ( .A0(n4009), .A1(n4010), .S(n1988), .Z(n4011) );
  CMXI2XL U2324 ( .A0(n1663), .A1(n1664), .S(net87791), .Z(n4997) );
  CMXI2XL U2325 ( .A0(n4275), .A1(n4276), .S(net87702), .Z(n4292) );
  CMXI2XL U2326 ( .A0(n1665), .A1(n1666), .S(net87809), .Z(n3971) );
  CIVXL U2327 ( .A(inst_fetch[1]), .Z(n1667) );
  CMXI2XL U2328 ( .A0(\reg_mem[2][13] ), .A1(\reg_mem[10][13] ), .S(net87537), 
        .Z(net79482) );
  CMXI2XL U2329 ( .A0(n3710), .A1(n1535), .S(n2174), .Z(n3711) );
  CMXI2XL U2330 ( .A0(n4155), .A1(n4156), .S(net87703), .Z(n4172) );
  CMXI2X1 U2331 ( .A0(n4993), .A1(n4994), .S(net87699), .Z(n4995) );
  CMXI2XL U2332 ( .A0(n1670), .A1(n1671), .S(net87807), .Z(n4834) );
  CMXI2X1 U2333 ( .A0(n4199), .A1(n4200), .S(net87703), .Z(n4216) );
  CIVXL U2334 ( .A(N118), .Z(n2789) );
  CMXI2XL U2335 ( .A0(n1672), .A1(n1673), .S(net87802), .Z(n3997) );
  CMXI2XL U2336 ( .A0(n1674), .A1(n1675), .S(net87804), .Z(n3998) );
  CMXI2X1 U2337 ( .A0(n3096), .A1(n3095), .S(n1450), .Z(n3097) );
  CMXI2X1 U2338 ( .A0(n2895), .A1(n2896), .S(net87483), .Z(n2897) );
  CMXI2X1 U2339 ( .A0(n3781), .A1(n3782), .S(net87697), .Z(n3798) );
  CMXI2XL U2340 ( .A0(n1676), .A1(n1677), .S(net87798), .Z(n4256) );
  CND2IXL U2341 ( .B(n2786), .A(n2785), .Z(alu_op_c[23]) );
  CMXI2XL U2342 ( .A0(n1678), .A1(n1679), .S(net87797), .Z(n5030) );
  CMXI2X1 U2343 ( .A0(n4455), .A1(n4456), .S(net87701), .Z(n4472) );
  CMXI2XL U2344 ( .A0(\reg_mem[1][13] ), .A1(\reg_mem[9][13] ), .S(net87519), 
        .Z(net79475) );
  CMXI2XL U2345 ( .A0(\reg_mem[0][13] ), .A1(\reg_mem[8][13] ), .S(net87542), 
        .Z(net79481) );
  CMXI2XL U2346 ( .A0(n1680), .A1(n1681), .S(net87800), .Z(n4002) );
  CMXI2X1 U2347 ( .A0(n4014), .A1(n4013), .S(net82865), .Z(n4040) );
  CMXI2X1 U2348 ( .A0(n4255), .A1(n4256), .S(n1988), .Z(n4257) );
  CMXI2XL U2349 ( .A0(\reg_mem[0][16] ), .A1(\reg_mem[1][16] ), .S(net87807), 
        .Z(n1682) );
  CMXI2XL U2350 ( .A0(\reg_mem[2][16] ), .A1(\reg_mem[3][16] ), .S(net87791), 
        .Z(n1683) );
  CANR4CX1 U2351 ( .A(n339), .B(n5241), .C(n5263), .D(opcode_ex[3]), .Z(n338)
         );
  CIVXL U2352 ( .A(n340), .Z(n5263) );
  CND2X1 U2353 ( .A(n2455), .B(i_type), .Z(n2040) );
  CMXI2XL U2354 ( .A0(net78600), .A1(net78599), .S(net87990), .Z(N230) );
  CMXI2XL U2355 ( .A0(net78476), .A1(net78475), .S(net87990), .Z(N228) );
  CIVX2 U2356 ( .A(n1684), .Z(n1686) );
  CNIVX1 U2357 ( .A(n1688), .Z(n1687) );
  CNIVX1 U2358 ( .A(prog_count_de[3]), .Z(n1688) );
  CNIVX1 U2359 ( .A(n1690), .Z(n1689) );
  CNIVX1 U2360 ( .A(prog_count_de[2]), .Z(n1690) );
  CAOR2X2 U2361 ( .A(\reg_mem[11][29] ), .B(n2304), .C(n2308), .D(n161), .Z(
        n994) );
  CIVDX1 U2362 ( .A(i_type), .Z1(n1692) );
  CIVDX1 U2363 ( .A(j_type), .Z1(n1695) );
  CNIVX1 U2364 ( .A(n1695), .Z(n1694) );
  CNIVX1 U2365 ( .A(n1697), .Z(n1696) );
  CNIVX1 U2366 ( .A(n1698), .Z(n1697) );
  CNIVX1 U2367 ( .A(regB[31]), .Z(n1698) );
  CIVXL U2368 ( .A(regB[29]), .Z(n1700) );
  CIVX2 U2369 ( .A(n1700), .Z(n1701) );
  CNIVX1 U2370 ( .A(n1703), .Z(n1702) );
  CNIVX1 U2371 ( .A(n1704), .Z(n1703) );
  CNIVX1 U2372 ( .A(regB[28]), .Z(n1704) );
  CNIVX1 U2373 ( .A(n1706), .Z(n1705) );
  CNIVX1 U2374 ( .A(n1707), .Z(n1706) );
  CNIVX1 U2375 ( .A(regB[27]), .Z(n1707) );
  CNIVX1 U2376 ( .A(n1709), .Z(n1708) );
  CNIVX1 U2377 ( .A(n1710), .Z(n1709) );
  CNIVX1 U2378 ( .A(regB[26]), .Z(n1710) );
  CNIVX1 U2379 ( .A(n1712), .Z(n1711) );
  CNIVX1 U2380 ( .A(n1713), .Z(n1712) );
  CNIVX1 U2381 ( .A(regB[25]), .Z(n1713) );
  CNIVX1 U2382 ( .A(n1715), .Z(n1714) );
  CNIVX1 U2383 ( .A(n1716), .Z(n1715) );
  CNIVX1 U2384 ( .A(regB[24]), .Z(n1716) );
  CNIVX1 U2385 ( .A(n2021), .Z(n1717) );
  CNIVX1 U2386 ( .A(n1719), .Z(n1718) );
  CNIVX1 U2387 ( .A(n1720), .Z(n1719) );
  CNIVX1 U2388 ( .A(regB[22]), .Z(n1720) );
  CNIVX1 U2389 ( .A(n1722), .Z(n1721) );
  CNIVX1 U2390 ( .A(n1723), .Z(n1722) );
  CNIVX1 U2391 ( .A(regB[21]), .Z(n1723) );
  CNIVX1 U2392 ( .A(n1725), .Z(n1724) );
  CNIVX1 U2393 ( .A(n1726), .Z(n1725) );
  CNIVX1 U2394 ( .A(regB[20]), .Z(n1726) );
  CNIVX1 U2395 ( .A(n1728), .Z(n1727) );
  CNIVX1 U2396 ( .A(n1729), .Z(n1728) );
  CNIVX1 U2397 ( .A(regB[19]), .Z(n1729) );
  CNIVX1 U2398 ( .A(n1731), .Z(n1730) );
  CNIVX1 U2399 ( .A(n2051), .Z(n1731) );
  CNIVX1 U2400 ( .A(n1733), .Z(n1732) );
  CNIVX1 U2401 ( .A(n2106), .Z(n1733) );
  CNIVX1 U2402 ( .A(n1735), .Z(n1734) );
  CNIVX1 U2403 ( .A(n1736), .Z(n1735) );
  CNIVX1 U2404 ( .A(regB[15]), .Z(n1736) );
  CIVX3 U2405 ( .A(n1737), .Z(n1738) );
  CIVXL U2406 ( .A(regB[14]), .Z(n1737) );
  CNIVX1 U2407 ( .A(n1740), .Z(n1739) );
  CNIVX1 U2408 ( .A(n1741), .Z(n1740) );
  CNIVX1 U2409 ( .A(n2026), .Z(n1741) );
  CNIVX1 U2410 ( .A(n1743), .Z(n1742) );
  CNIVX1 U2411 ( .A(n1744), .Z(n1743) );
  CNIVX1 U2412 ( .A(regB[12]), .Z(n1744) );
  CNIVX1 U2413 ( .A(n1746), .Z(n1745) );
  CNIVX1 U2414 ( .A(n2033), .Z(n1746) );
  CNIVX1 U2415 ( .A(n1748), .Z(n1747) );
  CNIVX1 U2416 ( .A(n1749), .Z(n1748) );
  CNIVX1 U2417 ( .A(regB[10]), .Z(n1749) );
  CNIVX1 U2418 ( .A(n1751), .Z(n1750) );
  CNIVX1 U2419 ( .A(n1752), .Z(n1751) );
  CNIVX1 U2420 ( .A(regB[9]), .Z(n1752) );
  CNIVX1 U2421 ( .A(n1754), .Z(n1753) );
  CNIVX1 U2422 ( .A(n1755), .Z(n1754) );
  CNIVX1 U2423 ( .A(regB[8]), .Z(n1755) );
  CNIVX1 U2424 ( .A(n1757), .Z(n1756) );
  CNIVX1 U2425 ( .A(n1758), .Z(n1757) );
  CNIVX1 U2426 ( .A(regB[7]), .Z(n1758) );
  CNIVX1 U2427 ( .A(n1760), .Z(n1759) );
  CNIVX1 U2428 ( .A(n1761), .Z(n1760) );
  CNIVX1 U2429 ( .A(regB[6]), .Z(n1761) );
  CNIVX1 U2430 ( .A(n2050), .Z(n1762) );
  CNIVX1 U2431 ( .A(n1764), .Z(n1763) );
  CNIVX1 U2432 ( .A(n2110), .Z(n1764) );
  CNIVX1 U2433 ( .A(n1766), .Z(n1765) );
  CNIVX1 U2434 ( .A(n1767), .Z(n1766) );
  CNIVX1 U2435 ( .A(n1686), .Z(n1767) );
  CNIVX1 U2436 ( .A(n1769), .Z(n1768) );
  CNIVX1 U2437 ( .A(n2047), .Z(n1769) );
  CIVX3 U2438 ( .A(n1770), .Z(n1771) );
  CIVXL U2439 ( .A(regB[1]), .Z(n1770) );
  CNIVX1 U2440 ( .A(n1773), .Z(n1772) );
  CNIVX1 U2441 ( .A(n1774), .Z(n1773) );
  CNIVX1 U2442 ( .A(regB[0]), .Z(n1774) );
  CNIVX1 U2443 ( .A(n1776), .Z(n1775) );
  CNIVX1 U2444 ( .A(alu_op[8]), .Z(n1776) );
  CNIVX1 U2445 ( .A(n1778), .Z(n1777) );
  CNIVX1 U2446 ( .A(alu_op[31]), .Z(n1778) );
  CNIVX1 U2447 ( .A(n1780), .Z(n1779) );
  CNIVX1 U2448 ( .A(alu_op[1]), .Z(n1780) );
  CNIVX1 U2449 ( .A(n1782), .Z(n1781) );
  CNIVX1 U2450 ( .A(alu_op[2]), .Z(n1782) );
  CNIVX1 U2451 ( .A(n1784), .Z(n1783) );
  CNIVX1 U2452 ( .A(alu_op[3]), .Z(n1784) );
  CNIVX1 U2453 ( .A(n1786), .Z(n1785) );
  CNIVX1 U2454 ( .A(alu_op[4]), .Z(n1786) );
  CNIVX1 U2455 ( .A(n1788), .Z(n1787) );
  CNIVX1 U2456 ( .A(alu_op[5]), .Z(n1788) );
  CNIVX1 U2457 ( .A(n1790), .Z(n1789) );
  CNIVX1 U2458 ( .A(alu_op[6]), .Z(n1790) );
  CNIVX1 U2459 ( .A(n1792), .Z(n1791) );
  CNIVX1 U2460 ( .A(alu_op[7]), .Z(n1792) );
  CNIVX1 U2461 ( .A(n1794), .Z(n1793) );
  CNIVX1 U2462 ( .A(alu_op[9]), .Z(n1794) );
  CNIVX1 U2463 ( .A(n1796), .Z(n1795) );
  CNIVX1 U2464 ( .A(alu_op[10]), .Z(n1796) );
  CNIVX1 U2465 ( .A(n1798), .Z(n1797) );
  CNIVX1 U2466 ( .A(alu_op[11]), .Z(n1798) );
  CNIVX1 U2467 ( .A(n1800), .Z(n1799) );
  CNIVX1 U2468 ( .A(alu_op[12]), .Z(n1800) );
  CNIVX1 U2469 ( .A(n1802), .Z(n1801) );
  CNIVX1 U2470 ( .A(alu_op[0]), .Z(n1802) );
  CNIVX1 U2471 ( .A(n1804), .Z(n1803) );
  CNIVX1 U2472 ( .A(alu_op[30]), .Z(n1804) );
  CNIVX1 U2473 ( .A(n1806), .Z(n1805) );
  CNIVX1 U2474 ( .A(alu_op[13]), .Z(n1806) );
  CNIVX1 U2475 ( .A(n1808), .Z(n1807) );
  CNIVX1 U2476 ( .A(alu_op[14]), .Z(n1808) );
  CNIVX1 U2477 ( .A(n1810), .Z(n1809) );
  CNIVX1 U2478 ( .A(alu_op[15]), .Z(n1810) );
  CNIVX1 U2479 ( .A(n1812), .Z(n1811) );
  CNIVX1 U2480 ( .A(alu_op[16]), .Z(n1812) );
  CNIVX1 U2481 ( .A(n1814), .Z(n1813) );
  CNIVX1 U2482 ( .A(alu_op[17]), .Z(n1814) );
  CNIVX1 U2483 ( .A(n1816), .Z(n1815) );
  CNIVX1 U2484 ( .A(alu_op[18]), .Z(n1816) );
  CNIVX1 U2485 ( .A(n1818), .Z(n1817) );
  CNIVX1 U2486 ( .A(alu_op[19]), .Z(n1818) );
  CNIVX1 U2487 ( .A(n1820), .Z(n1819) );
  CNIVX1 U2488 ( .A(alu_op[20]), .Z(n1820) );
  CNIVX1 U2489 ( .A(n1822), .Z(n1821) );
  CNIVX1 U2490 ( .A(alu_op[21]), .Z(n1822) );
  CNIVX1 U2491 ( .A(n1824), .Z(n1823) );
  CNIVX1 U2492 ( .A(alu_op[22]), .Z(n1824) );
  CNIVX1 U2493 ( .A(n1826), .Z(n1825) );
  CNIVX1 U2494 ( .A(alu_op[23]), .Z(n1826) );
  CNIVX1 U2495 ( .A(n1828), .Z(n1827) );
  CNIVX1 U2496 ( .A(alu_op[24]), .Z(n1828) );
  CNIVX1 U2497 ( .A(n1830), .Z(n1829) );
  CNIVX1 U2498 ( .A(alu_op[25]), .Z(n1830) );
  CNIVX1 U2499 ( .A(n1832), .Z(n1831) );
  CNIVX1 U2500 ( .A(alu_op[26]), .Z(n1832) );
  CNIVX1 U2501 ( .A(n1834), .Z(n1833) );
  CNIVX1 U2502 ( .A(alu_op[27]), .Z(n1834) );
  CNIVX1 U2503 ( .A(n1836), .Z(n1835) );
  CNIVX1 U2504 ( .A(alu_op[28]), .Z(n1836) );
  CNIVX1 U2505 ( .A(n1838), .Z(n1837) );
  CNIVX1 U2506 ( .A(alu_op[29]), .Z(n1838) );
  CNIVX1 U2507 ( .A(opcode_ex[5]), .Z(n1839) );
  CNIVX1 U2508 ( .A(opcode_ex[2]), .Z(n1840) );
  CNIVX1 U2509 ( .A(opcode_ex[4]), .Z(n1841) );
  CNIVX1 U2510 ( .A(opcode_ex[3]), .Z(n1842) );
  CAOR2X2 U2511 ( .A(\reg_mem[3][8] ), .B(net82537), .C(net82571), .D(n2226), 
        .Z(n1271) );
  CNIVX1 U2512 ( .A(opcode_ex[0]), .Z(n1843) );
  CDLY1XL U2513 ( .A(opcode_ex[1]), .Z(n1844) );
  CNIVX1 U2514 ( .A(n1846), .Z(n1845) );
  CNIVX1 U2515 ( .A(r_type_mem), .Z(n1846) );
  CIVDX1 U2516 ( .A(regc_addr_mem[4]), .Z1(n1849) );
  CNIVX1 U2517 ( .A(n1849), .Z(n1848) );
  CIVDX1 U2518 ( .A(regc_addr_mem[3]), .Z1(n1852) );
  CNIVX1 U2519 ( .A(n1852), .Z(n1851) );
  CIVDX1 U2520 ( .A(regc_addr_mem[1]), .Z1(n1855) );
  CNIVX1 U2521 ( .A(n1855), .Z(n1854) );
  CIVDX1 U2522 ( .A(regc_addr_mem[0]), .Z1(n1858) );
  CNIVX1 U2523 ( .A(n1858), .Z(n1857) );
  CIVDX1 U2524 ( .A(regc_addr_mem[2]), .Z1(n1861) );
  CNIVX1 U2525 ( .A(n1861), .Z(n1860) );
  CIVDX1 U2526 ( .A(regb_addr_mem[4]), .Z1(n1864) );
  CNIVX1 U2527 ( .A(n1864), .Z(n1863) );
  CIVDX1 U2528 ( .A(regb_addr_mem[3]), .Z1(n1867) );
  CNIVX1 U2529 ( .A(n1867), .Z(n1866) );
  CIVDX1 U2530 ( .A(regb_addr_mem[0]), .Z1(n1870) );
  CNIVX1 U2531 ( .A(n1870), .Z(n1869) );
  CIVDX1 U2532 ( .A(regb_addr_mem[2]), .Z1(n1873) );
  CNIVX1 U2533 ( .A(n1873), .Z(n1872) );
  CIVDX1 U2534 ( .A(regb_addr_mem[1]), .Z1(n1876) );
  CNIVX1 U2535 ( .A(n1876), .Z(n1875) );
  CNIVX1 U2536 ( .A(n1239), .Z(n1877) );
  CAOR2XL U2537 ( .A(\reg_mem[4][8] ), .B(net82497), .C(net82505), .D(n2227), 
        .Z(n1239) );
  CAOR2X2 U2538 ( .A(\reg_mem[5][8] ), .B(net82457), .C(net82491), .D(n182), 
        .Z(n1207) );
  CANR2XL U2539 ( .A(alu_op_c[3]), .B(n3750), .C(regA[3]), .D(n3739), .Z(n3487) );
  CIVDX1 U2540 ( .A(prog_count_de[7]), .Z1(n1880) );
  CNIVX1 U2541 ( .A(n1880), .Z(n1879) );
  CNIVX1 U2542 ( .A(prog_count_c[4]), .Z(n1881) );
  CIVDX1 U2543 ( .A(prog_count_de[0]), .Z1(n1884) );
  CNIVX1 U2544 ( .A(n1884), .Z(n1883) );
  CIVDX1 U2545 ( .A(prog_count_de[4]), .Z1(n1887) );
  CNIVX1 U2546 ( .A(n1887), .Z(n1886) );
  CIVDX1 U2547 ( .A(prog_count_de[5]), .Z1(n1890) );
  CNIVX1 U2548 ( .A(n1890), .Z(n1889) );
  CNIVX1 U2549 ( .A(n1892), .Z(n1891) );
  CNIVX1 U2550 ( .A(prog_count_de[1]), .Z(n1892) );
  CIVDX1 U2551 ( .A(prog_count_de[6]), .Z1(n1895) );
  CNIVX1 U2552 ( .A(n1895), .Z(n1894) );
  CNIVX1 U2553 ( .A(j_type_wb_c), .Z(n1896) );
  CAN3X4 U2554 ( .A(n243), .B(opcode_mem[2]), .C(i_type_mem), .Z(i_type_wb_c)
         );
  CIVDX1 U2555 ( .A(regc_addr[4]), .Z1(n1899) );
  CNIVX1 U2556 ( .A(n1899), .Z(n1898) );
  CIVDX1 U2557 ( .A(regc_addr[3]), .Z1(n1902) );
  CNIVX1 U2558 ( .A(n1902), .Z(n1901) );
  CIVDX1 U2559 ( .A(regc_addr[2]), .Z1(n1905) );
  CNIVX1 U2560 ( .A(n1905), .Z(n1904) );
  CIVDX1 U2561 ( .A(regc_addr[1]), .Z1(n1908) );
  CNIVX1 U2562 ( .A(n1908), .Z(n1907) );
  CIVDX1 U2563 ( .A(regc_addr[0]), .Z1(n1911) );
  CNIVX1 U2564 ( .A(n1911), .Z(n1910) );
  CIVDX1 U2565 ( .A(regb_addr[4]), .Z1(n1913) );
  CIVDX1 U2566 ( .A(regb_addr[3]), .Z1(n1915) );
  CIVDX1 U2567 ( .A(regb_addr[2]), .Z1(n1917) );
  CIVDX1 U2568 ( .A(regb_addr[1]), .Z1(n1919) );
  CNIVX1 U2569 ( .A(n1921), .Z(n1920) );
  CNIVX1 U2570 ( .A(regb_addr[0]), .Z(n1921) );
  CNIVX2 U2571 ( .A(N22), .Z(n1923) );
  CNIVX1 U2572 ( .A(n1923), .Z(n1922) );
  CNIVX1 U2573 ( .A(n1925), .Z(n1924) );
  CNIVX1 U2574 ( .A(prog_count_o[7]), .Z(n1925) );
  CIVDX1 U2575 ( .A(prog_count_o[4]), .Z1(n1927) );
  CIVDX1 U2576 ( .A(prog_count_o[5]), .Z1(n1929) );
  CNIVX2 U2577 ( .A(prog_count_o[6]), .Z(n1930) );
  CNIVX1 U2578 ( .A(r_type), .Z(n1931) );
  CNIVX2 U2579 ( .A(N23), .Z(n1933) );
  CNIVX1 U2580 ( .A(n1933), .Z(n1932) );
  CNIVX2 U2581 ( .A(prog_count_o[3]), .Z(n1935) );
  CIVX2 U2582 ( .A(n517), .Z(n1936) );
  CIVX2 U2583 ( .A(n1936), .Z(n1937) );
  CAOR2XL U2584 ( .A(\reg_mem[26][26] ), .B(n1501), .C(n1500), .D(n164), .Z(
        n517) );
  CNIVX2 U2585 ( .A(\reg_mem[20][29] ), .Z(n1938) );
  CAOR2XL U2586 ( .A(n1938), .B(n2351), .C(n2354), .D(n161), .Z(n706) );
  CNIVX1 U2587 ( .A(rst), .Z(n1939) );
  CNIVXL U2588 ( .A(n209), .Z(n1940) );
  CND3XL U2589 ( .A(n192), .B(n1939), .C(n210), .Z(n209) );
  CND2X1 U2590 ( .A(n1943), .B(n1944), .Z(n4985) );
  CIVX1 U2591 ( .A(n1988), .Z(n1945) );
  CND2X1 U2592 ( .A(n1947), .B(n1945), .Z(n1944) );
  CMXI2XL U2593 ( .A0(\reg_mem[4][27] ), .A1(\reg_mem[5][27] ), .S(net87800), 
        .Z(n1946) );
  CMXI2XL U2594 ( .A0(\reg_mem[6][27] ), .A1(\reg_mem[7][27] ), .S(net87802), 
        .Z(n1947) );
  CIVX1 U2595 ( .A(net86939), .Z(net87622) );
  CMXI2XL U2596 ( .A0(n1948), .A1(n1949), .S(net87794), .Z(n5034) );
  CMXI2X1 U2597 ( .A0(n4620), .A1(n4619), .S(net82863), .Z(n4646) );
  CMXI2XL U2598 ( .A0(n1950), .A1(n1951), .S(net87793), .Z(n4260) );
  CMXI2XL U2599 ( .A0(n1952), .A1(n1953), .S(net87797), .Z(net78626) );
  CMXI2XL U2600 ( .A0(n1954), .A1(n1955), .S(net87795), .Z(n4838) );
  CMXI2X1 U2601 ( .A0(n4171), .A1(n4172), .S(n1960), .Z(n4173) );
  CND2X1 U2602 ( .A(n1956), .B(n1957), .Z(n4608) );
  CND2XL U2603 ( .A(net87795), .B(\reg_mem[5][20] ), .Z(n1956) );
  CND2X1 U2604 ( .A(\reg_mem[4][20] ), .B(n1993), .Z(n1957) );
  CMXI2XL U2605 ( .A0(n1958), .A1(n1959), .S(net87802), .Z(n4251) );
  CMXI2X1 U2606 ( .A0(n3899), .A1(n3900), .S(n1988), .Z(n3901) );
  CMXI2X1 U2607 ( .A0(n3861), .A1(n3862), .S(n1960), .Z(net78599) );
  CMXI2X1 U2608 ( .A0(n4611), .A1(n4612), .S(n1988), .Z(n4618) );
  CNIVX3 U2609 ( .A(net87620), .Z(net87631) );
  CANR1X1 U2610 ( .A(N158), .B(n3701), .C(n2829), .Z(n2831) );
  CNR2IX1 U2611 ( .B(N117), .A(n2272), .Z(n2829) );
  CMXI2X1 U2612 ( .A0(n2511), .A1(n2512), .S(net87233), .Z(n2520) );
  CMXI2X1 U2613 ( .A0(n4149), .A1(n4150), .S(n1988), .Z(n4156) );
  CMXI2X1 U2614 ( .A0(n4268), .A1(n4267), .S(net82863), .Z(n4294) );
  CMXI2X1 U2615 ( .A0(n2687), .A1(n2688), .S(n1470), .Z(n2692) );
  CMXI2X1 U2616 ( .A0(n4861), .A1(n4891), .S(n2089), .Z(n2687) );
  CMXI2XL U2617 ( .A0(n1961), .A1(n1962), .S(net87809), .Z(n4095) );
  CMXI2XL U2618 ( .A0(n4517), .A1(n4518), .S(net87990), .Z(N215) );
  CMXI2XL U2619 ( .A0(net78041), .A1(net78042), .S(net86657), .Z(N221) );
  CIVDX1 U2620 ( .A(net15031), .Z0(n1960), .Z1(net82865) );
  CMXI2XL U2621 ( .A0(n1963), .A1(n1964), .S(net87797), .Z(n4493) );
  CMXI2X1 U2622 ( .A0(n4473), .A1(n4474), .S(net87990), .Z(N216) );
  CMXI2X1 U2623 ( .A0(n4001), .A1(n4002), .S(n1988), .Z(n4003) );
  CMXI2XL U2624 ( .A0(n1965), .A1(n1966), .S(net87804), .Z(n4005) );
  CMXI2X1 U2625 ( .A0(n2525), .A1(n2526), .S(net87233), .Z(n2534) );
  CMX2X1 U2626 ( .A0(\reg_mem[18][7] ), .A1(\reg_mem[19][7] ), .S(net87795), 
        .Z(n4059) );
  CMXI2X1 U2627 ( .A0(n3719), .A1(n3720), .S(net87508), .Z(n3736) );
  CND2X1 U2628 ( .A(n1967), .B(n1968), .Z(n4183) );
  CND2XL U2629 ( .A(net87795), .B(\reg_mem[11][10] ), .Z(n1967) );
  CND2X1 U2630 ( .A(\reg_mem[10][10] ), .B(n1993), .Z(n1968) );
  CAN2X1 U2631 ( .A(net87252), .B(net87538), .Z(n2142) );
  CMXI2XL U2632 ( .A0(n1969), .A1(n1970), .S(net87807), .Z(n4252) );
  CMXI2X1 U2633 ( .A0(n4601), .A1(n4602), .S(net87990), .Z(N213) );
  CMXI2X1 U2634 ( .A0(n4483), .A1(n4484), .S(n1988), .Z(n4490) );
  CIVX1 U2635 ( .A(alu_op_c[11]), .Z(n3213) );
  CMXI2X1 U2636 ( .A0(n4855), .A1(n4856), .S(net88175), .Z(n4857) );
  CMXI2X1 U2637 ( .A0(n3797), .A1(n3798), .S(net88175), .Z(n3799) );
  CMXI2XL U2638 ( .A0(n1971), .A1(n1972), .S(net87806), .Z(n4984) );
  CMXI2X1 U2639 ( .A0(n4515), .A1(n4516), .S(net88175), .Z(n4517) );
  CMX2X1 U2640 ( .A0(alu_op_c[17]), .A1(n2151), .S(n1534), .Z(N286) );
  CMXI2XL U2641 ( .A0(n1973), .A1(n1974), .S(net87799), .Z(n2000) );
  CMXI2XL U2642 ( .A0(n2655), .A1(n2654), .S(n2189), .Z(n2658) );
  CMXI2X1 U2643 ( .A0(n2521), .A1(n2522), .S(n1470), .Z(n2526) );
  CMXI2XL U2644 ( .A0(\reg_mem[13][31] ), .A1(\reg_mem[29][31] ), .S(n2093), 
        .Z(n3655) );
  CNIVX4 U2645 ( .A(net87374), .Z(net87387) );
  CMXI2X1 U2646 ( .A0(n4081), .A1(n4082), .S(net88175), .Z(n4083) );
  CMXI2XL U2647 ( .A0(n4130), .A1(n4129), .S(net86657), .Z(N224) );
  CMXI2X1 U2648 ( .A0(n4833), .A1(n4834), .S(n1988), .Z(n4840) );
  CMXI2X1 U2649 ( .A0(n3917), .A1(n3918), .S(net88175), .Z(n3919) );
  CMX2X1 U2650 ( .A0(n1977), .A1(n1978), .S(net87638), .Z(n5082) );
  CMXI2XL U2651 ( .A0(\reg_mem[8][29] ), .A1(\reg_mem[9][29] ), .S(net87797), 
        .Z(n1977) );
  CMXI2XL U2652 ( .A0(\reg_mem[10][29] ), .A1(\reg_mem[11][29] ), .S(net87803), 
        .Z(n1978) );
  CMXI2XL U2653 ( .A0(n3919), .A1(n3920), .S(net87990), .Z(N229) );
  CNIVX4 U2654 ( .A(net87376), .Z(net87396) );
  CMXI2XL U2655 ( .A0(n4646), .A1(n4645), .S(net86657), .Z(N212) );
  CMXI2X1 U2656 ( .A0(n2724), .A1(n2725), .S(n2173), .Z(n2729) );
  CMXI2XL U2657 ( .A0(n4936), .A1(n4966), .S(n2081), .Z(n2655) );
  CMXI2XL U2658 ( .A0(\reg_mem[5][20] ), .A1(\reg_mem[13][20] ), .S(net87537), 
        .Z(n2879) );
  CMX2X1 U2659 ( .A0(n1979), .A1(n1980), .S(net87627), .Z(n4576) );
  CMXI2XL U2660 ( .A0(\reg_mem[8][19] ), .A1(\reg_mem[9][19] ), .S(net87803), 
        .Z(n1979) );
  CMXI2XL U2661 ( .A0(\reg_mem[10][19] ), .A1(\reg_mem[11][19] ), .S(net87803), 
        .Z(n1980) );
  CMXI2XL U2662 ( .A0(n4173), .A1(n4174), .S(net87990), .Z(N223) );
  CMXI2X1 U2663 ( .A0(n4983), .A1(n4984), .S(n1988), .Z(n4986) );
  CMXI2XL U2664 ( .A0(n4718), .A1(n4732), .S(net87544), .Z(n2800) );
  CMXI2X1 U2665 ( .A0(\reg_mem[4][29] ), .A1(\reg_mem[20][29] ), .S(n2090), 
        .Z(n2510) );
  CNIVX3 U2666 ( .A(n2079), .Z(n2090) );
  CMXI2XL U2667 ( .A0(n3799), .A1(n3800), .S(net87990), .Z(N232) );
  CMXI2XL U2668 ( .A0(n4294), .A1(n4293), .S(net86657), .Z(N220) );
  CMXI2XL U2669 ( .A0(n4938), .A1(n4968), .S(n2096), .Z(n2654) );
  CMXI2X1 U2670 ( .A0(n2947), .A1(n2948), .S(n2173), .Z(n2949) );
  CND2X1 U2671 ( .A(n1986), .B(n1987), .Z(net78090) );
  CND2X1 U2672 ( .A(n1990), .B(n1988), .Z(n1987) );
  CMXI2XL U2673 ( .A0(\reg_mem[6][11] ), .A1(\reg_mem[7][11] ), .S(net87799), 
        .Z(n1989) );
  CMXI2XL U2674 ( .A0(\reg_mem[4][11] ), .A1(\reg_mem[5][11] ), .S(net87799), 
        .Z(n1990) );
  CND2X1 U2675 ( .A(n1991), .B(n1992), .Z(n2004) );
  CND2XL U2676 ( .A(net87799), .B(\reg_mem[17][2] ), .Z(n1991) );
  CND2X1 U2677 ( .A(\reg_mem[16][2] ), .B(n1993), .Z(n1992) );
  CNIVX3 U2678 ( .A(net87514), .Z(net87530) );
  CND2X1 U2679 ( .A(n1994), .B(n1995), .Z(n2005) );
  CND2XL U2680 ( .A(net87799), .B(\reg_mem[17][4] ), .Z(n1994) );
  CND2X1 U2681 ( .A(\reg_mem[16][4] ), .B(n1993), .Z(n1995) );
  CIVX2 U2682 ( .A(inst_fetch[22]), .Z(n2001) );
  CNIVX8 U2683 ( .A(net87786), .Z(net87799) );
  CNIVX8 U2684 ( .A(net87789), .Z(net87800) );
  CNIVX8 U2685 ( .A(net87787), .Z(net87798) );
  CNR2IX1 U2686 ( .B(inst_fetch[22]), .A(net76768), .Z(net76777) );
  CMXI2X1 U2687 ( .A0(net77950), .A1(net77949), .S(net88175), .Z(net77917) );
  CMXI2XL U2688 ( .A0(net77918), .A1(net77917), .S(net87990), .Z(N219) );
  CIVDX1 U2689 ( .A(net15031), .Z0(net88175), .Z1(net82863) );
  CMXI2X1 U2690 ( .A0(net78478), .A1(net78477), .S(net88175), .Z(net78476) );
  CMXI2X1 U2691 ( .A0(net78602), .A1(net78601), .S(net88175), .Z(net78600) );
  CIVX2 U2692 ( .A(net78759), .Z(net15031) );
  CMXI2X1 U2693 ( .A0(net77966), .A1(net77965), .S(net87701), .Z(net77949) );
  CIVX1 U2694 ( .A(net86659), .Z(net87701) );
  CNIVX3 U2695 ( .A(net87622), .Z(net87638) );
  CNIVX3 U2696 ( .A(net87622), .Z(net87636) );
  CNIVX3 U2697 ( .A(net87622), .Z(net87635) );
  CNIVX8 U2698 ( .A(net87788), .Z(net87795) );
  CNIVX8 U2699 ( .A(net87786), .Z(net87797) );
  CNIVX8 U2700 ( .A(net87789), .Z(net87794) );
  CMXI2X1 U2701 ( .A0(net77967), .A1(n2002), .S(net87636), .Z(net77966) );
  CMXI2X1 U2702 ( .A0(net77969), .A1(net77970), .S(net87802), .Z(n2002) );
  CNIVX8 U2703 ( .A(net87788), .Z(net87803) );
  CNIVX8 U2704 ( .A(net87787), .Z(net87804) );
  CND2IXL U2705 ( .B(n2003), .A(net87488), .Z(net86939) );
  CIVX2 U2706 ( .A(inst_fetch[23]), .Z(n2003) );
  CMXI2X1 U2707 ( .A0(\reg_mem[3][13] ), .A1(\reg_mem[11][13] ), .S(net87532), 
        .Z(net79476) );
  CNR2IX1 U2708 ( .B(inst_fetch[23]), .A(net76768), .Z(net76776) );
  CNIVX8 U2709 ( .A(net87789), .Z(net87802) );
  CIVX2 U2710 ( .A(\reg_mem[7][13] ), .Z(net77970) );
  CIVX2 U2711 ( .A(\reg_mem[6][13] ), .Z(net77969) );
  CMXI2X1 U2712 ( .A0(\reg_mem[0][11] ), .A1(\reg_mem[4][11] ), .S(net87258), 
        .Z(net79408) );
  CMXI2X1 U2713 ( .A0(\reg_mem[1][11] ), .A1(\reg_mem[5][11] ), .S(net87277), 
        .Z(net79406) );
  CMXI2X1 U2714 ( .A0(net78089), .A1(net78090), .S(net87717), .Z(net78073) );
  CIVX1 U2715 ( .A(net87700), .Z(net87717) );
  CIVXL U2716 ( .A(net86659), .Z(net87700) );
  CIVX1 U2717 ( .A(net87700), .Z(net87719) );
  CIVX1 U2718 ( .A(net87700), .Z(net87718) );
  CIVX1 U2719 ( .A(net87700), .Z(net87716) );
  CNIVX3 U2720 ( .A(net87622), .Z(net87642) );
  CNIVX3 U2721 ( .A(net87622), .Z(net87640) );
  CNIVX3 U2722 ( .A(net87622), .Z(net87639) );
  CMXI2X1 U2723 ( .A0(net78097), .A1(net78098), .S(net87634), .Z(net78089) );
  CNIVX3 U2724 ( .A(net87620), .Z(net87634) );
  CIVXL U2725 ( .A(net86939), .Z(net87620) );
  CMXI2X1 U2726 ( .A0(\reg_mem[3][11] ), .A1(\reg_mem[7][11] ), .S(net87263), 
        .Z(net79407) );
  CMXI2X1 U2727 ( .A0(\reg_mem[2][11] ), .A1(\reg_mem[6][11] ), .S(net87248), 
        .Z(net79409) );
  CNIVX3 U2728 ( .A(net87620), .Z(net87633) );
  CNIVX3 U2729 ( .A(net87620), .Z(net87632) );
  CMX2XL U2730 ( .A0(\reg_mem[2][11] ), .A1(\reg_mem[3][11] ), .S(net87790), 
        .Z(net78098) );
  CMXI2X1 U2731 ( .A0(n2004), .A1(net78626), .S(net87625), .Z(net78617) );
  CMXI2X1 U2732 ( .A0(\reg_mem[16][2] ), .A1(\reg_mem[17][2] ), .S(net87409), 
        .Z(net79032) );
  CMXI2X1 U2733 ( .A0(net78618), .A1(net78617), .S(net87701), .Z(net78601) );
  CNIVX3 U2734 ( .A(net87618), .Z(net87625) );
  CIVXL U2735 ( .A(net86939), .Z(net87618) );
  CNIVX3 U2736 ( .A(net87618), .Z(net87626) );
  CNIVX3 U2737 ( .A(net87618), .Z(net87624) );
  CMXI2X1 U2738 ( .A0(net78619), .A1(net78620), .S(net87642), .Z(net78618) );
  CMXI2XL U2739 ( .A0(\reg_mem[18][2] ), .A1(\reg_mem[19][2] ), .S(net87407), 
        .Z(net79033) );
  CMXI2X1 U2740 ( .A0(net78621), .A1(net78622), .S(net87793), .Z(net78620) );
  CNIVX8 U2741 ( .A(net87786), .Z(net87793) );
  CNIVX8 U2742 ( .A(net87786), .Z(net87791) );
  CMXI2X1 U2743 ( .A0(n2005), .A1(net78502), .S(net87642), .Z(net78493) );
  CMXI2X1 U2744 ( .A0(\reg_mem[16][4] ), .A1(\reg_mem[17][4] ), .S(net87405), 
        .Z(net79122) );
  CMXI2X1 U2745 ( .A0(net78494), .A1(net78493), .S(net87701), .Z(net78477) );
  CND3X2 U2746 ( .A(net80175), .B(net76798), .C(net80176), .Z(net87488) );
  CANR1X2 U2747 ( .A(net80185), .B(net78795), .C(net80186), .Z(net80175) );
  CND3X2 U2748 ( .A(net80175), .B(net80176), .C(net76798), .Z(net78726) );
  CND3X1 U2749 ( .A(net80175), .B(net76798), .C(net80176), .Z(net87489) );
  CNR2X2 U2750 ( .A(n2008), .B(net78798), .Z(net80186) );
  CND3X1 U2751 ( .A(net78797), .B(inst_fetch[2]), .C(n2011), .Z(n2008) );
  CIVXL U2752 ( .A(inst_fetch[5]), .Z(n2011) );
  CIVXL U2753 ( .A(n2011), .Z(net87691) );
  CNR2X1 U2754 ( .A(n2009), .B(n2010), .Z(net80185) );
  CIVXL U2755 ( .A(n2012), .Z(n2010) );
  CIVXL U2756 ( .A(inst_fetch[5]), .Z(n2012) );
  CND2XL U2757 ( .A(inst_fetch[2]), .B(inst_fetch[4]), .Z(n2009) );
  CND2X2 U2758 ( .A(net80177), .B(net80178), .Z(net76798) );
  CND3X1 U2759 ( .A(n2006), .B(n2007), .C(net86647), .Z(net80176) );
  CNR2XL U2760 ( .A(inst_fetch[0]), .B(inst_fetch[4]), .Z(n2007) );
  CNR2XL U2761 ( .A(inst_fetch[3]), .B(n2012), .Z(n2006) );
  COND4CXL U2762 ( .A(inst_fetch[4]), .B(net78795), .C(net86675), .D(net88116), 
        .Z(net78792) );
  CIVXL U2763 ( .A(net78798), .Z(net78793) );
  CAN2XL U2764 ( .A(inst_fetch[5]), .B(inst_fetch[4]), .Z(net83592) );
  CAN2XL U2765 ( .A(inst_fetch[0]), .B(inst_fetch[1]), .Z(net86999) );
  CAN2XL U2766 ( .A(inst_fetch[2]), .B(inst_fetch[1]), .Z(net86647) );
  CND2XL U2767 ( .A(net80177), .B(n1479), .Z(net88101) );
  CND2XL U2768 ( .A(net78793), .B(net86647), .Z(net76796) );
  CMXI2X1 U2769 ( .A0(\reg_mem[18][4] ), .A1(\reg_mem[19][4] ), .S(net87411), 
        .Z(net79123) );
  CMXI2X1 U2770 ( .A0(net78497), .A1(net78498), .S(net87803), .Z(net78496) );
  CMXI2X1 U2771 ( .A0(net87836), .A1(n1667), .S(net87781), .Z(net78795) );
  CIVX1 U2772 ( .A(inst_fetch[0]), .Z(net87781) );
  CIVX1 U2773 ( .A(net87781), .Z(net87782) );
  CIVXL U2774 ( .A(net87835), .Z(net87836) );
  CIVXL U2775 ( .A(inst_fetch[3]), .Z(net87835) );
  CNR2X1 U2776 ( .A(inst_fetch[0]), .B(inst_fetch[4]), .Z(n2013) );
  CMXI2XL U2777 ( .A0(n4857), .A1(n4858), .S(net87990), .Z(N208) );
  CMXI2XL U2778 ( .A0(n4083), .A1(n4084), .S(net87990), .Z(N225) );
  CNIVX3 U2779 ( .A(n2078), .Z(n2104) );
  CMXI2X1 U2780 ( .A0(n2818), .A1(n1536), .S(n1471), .Z(n2819) );
  CMXI2X1 U2781 ( .A0(n2744), .A1(n2745), .S(net87508), .Z(n2746) );
  CMXI2X1 U2782 ( .A0(n2955), .A1(n2956), .S(net87233), .Z(n2957) );
  CIVX2 U2783 ( .A(n2014), .Z(n2016) );
  CMX2X1 U2784 ( .A0(n2017), .A1(n2018), .S(net87631), .Z(n5028) );
  CMXI2XL U2785 ( .A0(\reg_mem[0][28] ), .A1(\reg_mem[1][28] ), .S(net87790), 
        .Z(n2017) );
  CMXI2XL U2786 ( .A0(\reg_mem[2][28] ), .A1(\reg_mem[3][28] ), .S(net87803), 
        .Z(n2018) );
  CND2IX1 U2787 ( .B(net87483), .A(n2148), .Z(n3653) );
  CMXI2X1 U2788 ( .A0(n2644), .A1(n2645), .S(net87233), .Z(n2646) );
  CIVX1 U2789 ( .A(n2019), .Z(n2021) );
  CMXI2XL U2790 ( .A0(\reg_mem[15][31] ), .A1(\reg_mem[31][31] ), .S(n2090), 
        .Z(n3654) );
  CIVX2 U2791 ( .A(n2091), .Z(n2073) );
  CMXI2X1 U2792 ( .A0(n4481), .A1(n4482), .S(net87701), .Z(n4492) );
  CMXI2X1 U2793 ( .A0(n2969), .A1(n2970), .S(net87233), .Z(n2971) );
  CMXI2X1 U2794 ( .A0(\reg_mem[22][20] ), .A1(\reg_mem[30][20] ), .S(net87537), 
        .Z(n2886) );
  CMXI2X1 U2795 ( .A0(n4182), .A1(n4181), .S(net87727), .Z(n4192) );
  COND1X1 U2796 ( .A(n3604), .B(n2639), .C(n3615), .Z(n2663) );
  CMXI2X1 U2797 ( .A0(n3105), .A1(n3106), .S(net87233), .Z(n3114) );
  CMXI2X1 U2798 ( .A0(n3093), .A1(n3094), .S(n2173), .Z(n3098) );
  CIVX2 U2799 ( .A(n2023), .Z(n2025) );
  CMXI2XL U2800 ( .A0(n2155), .A1(n3742), .S(prog_count_o[6]), .Z(n3347) );
  CNIVX3 U2801 ( .A(n2077), .Z(n2103) );
  CMXI2X1 U2802 ( .A0(n3090), .A1(n3089), .S(n2200), .Z(n3091) );
  CMX2XL U2803 ( .A0(n2141), .A1(n3595), .S(n2114), .Z(N270) );
  CMXI2X1 U2804 ( .A0(n2727), .A1(n2726), .S(n2180), .Z(n2728) );
  CMXI2XL U2805 ( .A0(n3111), .A1(n3112), .S(net87233), .Z(n3113) );
  CMXI2X1 U2806 ( .A0(n4499), .A1(n4500), .S(net87701), .Z(n4516) );
  CMXI2XL U2807 ( .A0(\reg_mem[4][28] ), .A1(\reg_mem[20][28] ), .S(n2090), 
        .Z(n2556) );
  CIVX3 U2808 ( .A(n2173), .Z(n2200) );
  CIVXL U2809 ( .A(n3696), .Z(n3707) );
  COND3X1 U2810 ( .A(n2272), .B(n3391), .C(n3390), .D(n3389), .Z(alu_op_c[5])
         );
  CANR1X2 U2811 ( .A(N174), .B(n3704), .C(n3388), .Z(n3389) );
  CMXI2XL U2812 ( .A0(n2027), .A1(n2028), .S(net87799), .Z(n3858) );
  CMXI2XL U2813 ( .A0(n3578), .A1(n3577), .S(net87403), .Z(n3579) );
  CMXI2X1 U2814 ( .A0(n3857), .A1(n3858), .S(net88166), .Z(n3859) );
  CANR2XL U2815 ( .A(N188), .B(n3704), .C(N156), .D(n3701), .Z(n2909) );
  CIVXL U2816 ( .A(n1667), .Z(net88155) );
  CMXI2XL U2817 ( .A0(n4040), .A1(n4039), .S(net86657), .Z(N226) );
  CMXI2XL U2818 ( .A0(n2031), .A1(n2032), .S(net87799), .Z(n3854) );
  CMXI2X1 U2819 ( .A0(n2519), .A1(n2520), .S(net87508), .Z(n2536) );
  CIVX1 U2820 ( .A(n2069), .Z(n2067) );
  CMXI2X1 U2821 ( .A0(n4493), .A1(n4494), .S(n1988), .Z(n4500) );
  CMXI2XL U2822 ( .A0(n4814), .A1(n4813), .S(net86657), .Z(N209) );
  CIVXL U2823 ( .A(n1472), .Z(net87516) );
  CIVX2 U2824 ( .A(net83575), .Z(net87514) );
  CMXI2X1 U2825 ( .A0(n2657), .A1(n2658), .S(net87233), .Z(n2659) );
  COND1X1 U2826 ( .A(n2678), .B(n3604), .C(n3615), .Z(n2706) );
  CIVX3 U2827 ( .A(n2188), .Z(n2164) );
  CMXI2X1 U2828 ( .A0(n1457), .A1(n3557), .S(n1459), .Z(N271) );
  CMXI2X1 U2829 ( .A0(n3596), .A1(n2034), .S(n1534), .Z(n2141) );
  CMX2X1 U2830 ( .A0(n3580), .A1(n3579), .S(n1532), .Z(n2034) );
  CIVXL U2831 ( .A(inst_fetch[2]), .Z(net88115) );
  CIVX2 U2832 ( .A(net88115), .Z(net88116) );
  CIVX2 U2833 ( .A(n2035), .Z(n2037) );
  CIVX2 U2834 ( .A(n2167), .Z(n2038) );
  CIVX2 U2835 ( .A(n2167), .Z(n2039) );
  CIVX4 U2836 ( .A(n2461), .Z(n2167) );
  CNIVX3 U2837 ( .A(n2078), .Z(n2102) );
  CNIVX3 U2838 ( .A(n2076), .Z(n2101) );
  CNIVX3 U2839 ( .A(n2076), .Z(n2094) );
  CNIVX4 U2840 ( .A(n2079), .Z(n2080) );
  CMXI2XL U2841 ( .A0(\reg_mem[12][30] ), .A1(\reg_mem[28][30] ), .S(n2084), 
        .Z(n3619) );
  CMXI2XL U2842 ( .A0(\reg_mem[0][27] ), .A1(\reg_mem[16][27] ), .S(n2085), 
        .Z(n2596) );
  CIVX1 U2843 ( .A(net79756), .Z(net87380) );
  CMXI2X1 U2844 ( .A0(n2535), .A1(n2536), .S(net87483), .Z(n2537) );
  CIVX2 U2845 ( .A(n2118), .Z(n2119) );
  CIVX2 U2846 ( .A(n2040), .Z(n2041) );
  CANR1XL U2847 ( .A(n2454), .B(n2452), .C(n2451), .Z(n2042) );
  CIVX1 U2848 ( .A(n3344), .Z(n2456) );
  CMXI2XL U2849 ( .A0(n3145), .A1(n1468), .S(n2114), .Z(N282) );
  CND2IXL U2850 ( .B(n2717), .A(n2716), .Z(alu_op_c[24]) );
  CND2IX2 U2851 ( .B(n2043), .A(net78726), .Z(n2805) );
  CMXI2X1 U2852 ( .A0(\reg_mem[3][29] ), .A1(\reg_mem[19][29] ), .S(n1975), 
        .Z(n2521) );
  CMXI2XL U2853 ( .A0(n4562), .A1(n4561), .S(net86657), .Z(N214) );
  CMXI2X1 U2854 ( .A0(n3853), .A1(n3854), .S(n1988), .Z(n3860) );
  CMXI2X1 U2855 ( .A0(n4491), .A1(n4492), .S(net78759), .Z(n4518) );
  CMXI2XL U2856 ( .A0(n3995), .A1(n3996), .S(net87990), .Z(N227) );
  CAN2X4 U2857 ( .A(inst_fetch[26]), .B(n1478), .Z(net86657) );
  CMX2X1 U2858 ( .A0(n2044), .A1(n2045), .S(net87623), .Z(n4584) );
  CMXI2XL U2859 ( .A0(\reg_mem[16][19] ), .A1(\reg_mem[17][19] ), .S(net87797), 
        .Z(n2044) );
  CMXI2XL U2860 ( .A0(\reg_mem[18][19] ), .A1(\reg_mem[19][19] ), .S(net87790), 
        .Z(n2045) );
  CIVXL U2861 ( .A(immi_val[3]), .Z(n2046) );
  CND2XL U2862 ( .A(N184), .B(n3704), .Z(n3080) );
  CND2X1 U2863 ( .A(n2944), .B(n2943), .Z(alu_op_c[18]) );
  CND2X1 U2864 ( .A(n2814), .B(n1469), .Z(n2122) );
  CIVX2 U2865 ( .A(n2048), .Z(n2050) );
  CIVX1 U2866 ( .A(net79770), .Z(net87241) );
  CMX2X1 U2867 ( .A0(\reg_mem[1][22] ), .A1(\reg_mem[9][22] ), .S(net87523), 
        .Z(n2815) );
  CAN2X2 U2868 ( .A(net87488), .B(inst_fetch[27]), .Z(n2053) );
  CMXI2XL U2869 ( .A0(n2556), .A1(n2555), .S(n2184), .Z(n2557) );
  CMXI2XL U2870 ( .A0(n2836), .A1(n2835), .S(n2165), .Z(n2837) );
  CMXI2XL U2871 ( .A0(n3651), .A1(n3650), .S(n2183), .Z(n3652) );
  CMXI2XL U2872 ( .A0(n3029), .A1(n3028), .S(n2183), .Z(n3033) );
  CMXI2XL U2873 ( .A0(n2817), .A1(n2816), .S(n2183), .Z(n2818) );
  CMX2XL U2874 ( .A0(\reg_mem[16][17] ), .A1(\reg_mem[17][17] ), .S(net87790), 
        .Z(n4494) );
  CMX2XL U2875 ( .A0(\reg_mem[12][14] ), .A1(\reg_mem[13][14] ), .S(net87790), 
        .Z(n4340) );
  CMXI2X1 U2876 ( .A0(n2968), .A1(n2967), .S(n2198), .Z(n2969) );
  CMXI2X1 U2877 ( .A0(n3735), .A1(n3736), .S(n2075), .Z(n3738) );
  CNIVX4 U2878 ( .A(net87511), .Z(net87537) );
  CMXI2XL U2879 ( .A0(n3830), .A1(n3829), .S(net87795), .Z(n3831) );
  CMXI2XL U2880 ( .A0(n4210), .A1(n4209), .S(net87790), .Z(n4211) );
  CMXI2XL U2881 ( .A0(n4222), .A1(n4221), .S(net87809), .Z(n4223) );
  CMXI2XL U2882 ( .A0(n3982), .A1(n3981), .S(net87790), .Z(n3983) );
  CMXI2XL U2883 ( .A0(n5104), .A1(n5103), .S(net87806), .Z(n5108) );
  CMXI2XL U2884 ( .A0(n4836), .A1(n4835), .S(net87795), .Z(n4837) );
  CMXI2XL U2885 ( .A0(n4636), .A1(n4635), .S(net87797), .Z(n4640) );
  CMXI2XL U2886 ( .A0(n4624), .A1(n4623), .S(net87807), .Z(n4625) );
  CMXI2XL U2887 ( .A0(n5192), .A1(n5191), .S(net87804), .Z(n5193) );
  CMXI2XL U2888 ( .A0(n4880), .A1(n4879), .S(net87798), .Z(n4884) );
  CMXI2XL U2889 ( .A0(n4416), .A1(n4415), .S(net87795), .Z(n4420) );
  CMXI2XL U2890 ( .A0(n4868), .A1(n4867), .S(net87802), .Z(n4869) );
  CMXI2XL U2891 ( .A0(n4024), .A1(n4023), .S(net87802), .Z(n4028) );
  CMXI2XL U2892 ( .A0(n4402), .A1(n4401), .S(net87795), .Z(n4406) );
  CMX2XL U2893 ( .A0(\reg_mem[10][28] ), .A1(\reg_mem[11][28] ), .S(net87790), 
        .Z(n5029) );
  CMX2XL U2894 ( .A0(\reg_mem[8][30] ), .A1(\reg_mem[9][30] ), .S(net87790), 
        .Z(n5124) );
  CMX2XL U2895 ( .A0(\reg_mem[0][1] ), .A1(\reg_mem[1][1] ), .S(net87790), .Z(
        n3802) );
  CMX2XL U2896 ( .A0(\reg_mem[8][5] ), .A1(\reg_mem[9][5] ), .S(net87790), .Z(
        n3962) );
  CNR4X2 U2897 ( .A(n2706), .B(n2703), .C(n2704), .D(n2705), .Z(n2707) );
  CNR2IX1 U2898 ( .B(n2686), .A(n2685), .Z(n2705) );
  CND2XL U2899 ( .A(N191), .B(n3704), .Z(n2827) );
  COND1XL U2900 ( .A(n3563), .B(prog_count_o[5]), .C(n3343), .Z(n3742) );
  CAN3X2 U2901 ( .A(n3329), .B(n3330), .C(enable), .Z(n2153) );
  CMXI2X1 U2902 ( .A0(n3282), .A1(n3281), .S(n2096), .Z(n3284) );
  CIVX1 U2903 ( .A(net79756), .Z(net87378) );
  CNIVX2 U2904 ( .A(net87378), .Z(net87401) );
  CNIVX2 U2905 ( .A(net87378), .Z(net87404) );
  CMXI2X1 U2906 ( .A0(n3709), .A1(n3708), .S(n2200), .Z(n3712) );
  CND2X1 U2907 ( .A(n2746), .B(net87863), .Z(n2054) );
  CND2XL U2908 ( .A(n2747), .B(net87483), .Z(n2055) );
  CIVX2 U2909 ( .A(net87483), .Z(net87863) );
  CMX2XL U2910 ( .A0(alu_op_c[24]), .A1(n2149), .S(n1534), .Z(N293) );
  CIVX2 U2911 ( .A(n2056), .Z(n2058) );
  CNIVX8 U2912 ( .A(net87787), .Z(net87806) );
  CNIVX8 U2913 ( .A(net87787), .Z(net87807) );
  CNIVX8 U2914 ( .A(net87789), .Z(net87809) );
  CMXI2X1 U2915 ( .A0(n2721), .A1(n2720), .S(n1469), .Z(n2722) );
  CNIVX3 U2916 ( .A(n2078), .Z(n2100) );
  CNIVX3 U2917 ( .A(n2077), .Z(n2083) );
  CNIVX3 U2918 ( .A(n2079), .Z(n2084) );
  CMXI2X1 U2919 ( .A0(n2961), .A1(n2962), .S(n2175), .Z(n2963) );
  CMXI2X1 U2920 ( .A0(n2699), .A1(n2700), .S(net87233), .Z(n2701) );
  CIVXL U2921 ( .A(net86659), .Z(net87697) );
  CIVXL U2922 ( .A(net86659), .Z(net87698) );
  CIVXL U2923 ( .A(net86659), .Z(net87699) );
  CIVXL U2924 ( .A(net86659), .Z(net87702) );
  CIVXL U2925 ( .A(net86659), .Z(net87703) );
  CIVX1 U2926 ( .A(net87697), .Z(net87704) );
  CIVX1 U2927 ( .A(net87697), .Z(net87705) );
  CIVX1 U2928 ( .A(net87697), .Z(net87706) );
  CIVX1 U2929 ( .A(net87698), .Z(net87708) );
  CIVX1 U2930 ( .A(net87698), .Z(net87709) );
  CIVX1 U2931 ( .A(net87698), .Z(net87710) );
  CIVX1 U2932 ( .A(net87699), .Z(net87714) );
  CIVX1 U2933 ( .A(net87699), .Z(net87715) );
  CIVX1 U2934 ( .A(net87701), .Z(net87720) );
  CIVX1 U2935 ( .A(net87701), .Z(net87722) );
  CIVX1 U2936 ( .A(net87701), .Z(net87723) );
  CIVX1 U2937 ( .A(net87702), .Z(net87724) );
  CIVX1 U2938 ( .A(net87702), .Z(net87725) );
  CIVX1 U2939 ( .A(net87702), .Z(net87727) );
  CIVX1 U2940 ( .A(net87703), .Z(net87728) );
  CIVX1 U2941 ( .A(net87703), .Z(net87730) );
  CND2XL U2942 ( .A(N90), .B(n3697), .Z(n2631) );
  CND2IXL U2943 ( .B(n3698), .A(n3697), .Z(n3706) );
  CND2XL U2944 ( .A(N91), .B(n3697), .Z(n2622) );
  CND2XL U2945 ( .A(N92), .B(n3697), .Z(n2580) );
  CND2IXL U2946 ( .B(n3429), .A(n3697), .Z(n3435) );
  CND2XL U2947 ( .A(N94), .B(n3697), .Z(n3636) );
  CND2XL U2948 ( .A(N87), .B(n3697), .Z(n2781) );
  CND2XL U2949 ( .A(N85), .B(n3697), .Z(n2830) );
  CND2XL U2950 ( .A(N88), .B(n3697), .Z(n2714) );
  CND2IXL U2951 ( .B(n3040), .A(n3697), .Z(n3041) );
  CND2IXL U2952 ( .B(n3381), .A(n3697), .Z(n3390) );
  CND2XL U2953 ( .A(N86), .B(n3697), .Z(n2787) );
  CNIVX3 U2954 ( .A(n2076), .Z(n2099) );
  CMXI2X1 U2955 ( .A0(n3737), .A1(n3738), .S(n1534), .Z(N277) );
  CIVX2 U2956 ( .A(n2805), .Z(n2079) );
  CMXI2XL U2957 ( .A0(n2152), .A1(n2656), .S(n2176), .Z(n2657) );
  CMXI2X1 U2958 ( .A0(n4972), .A1(n4942), .S(n2073), .Z(n2152) );
  CND2X1 U2959 ( .A(N199), .B(n3704), .Z(n3642) );
  CIVX2 U2960 ( .A(n2061), .Z(n2062) );
  CIVXL U2961 ( .A(net87526), .Z(net87507) );
  CMX2X1 U2962 ( .A0(n4085), .A1(n4086), .S(n2066), .Z(n3709) );
  CND2X2 U2963 ( .A(net87489), .B(inst_fetch[29]), .Z(net79770) );
  CND2X2 U2964 ( .A(net87488), .B(inst_fetch[28]), .Z(n2461) );
  COND3XL U2965 ( .A(n2123), .B(n3084), .C(n3083), .D(n3082), .Z(n3086) );
  CNR2IXL U2966 ( .B(N106), .A(n2123), .Z(n3215) );
  CNR2IXL U2967 ( .B(N102), .A(n2272), .Z(n3326) );
  CIVXL U2968 ( .A(net86939), .Z(net87619) );
  CNIVX3 U2969 ( .A(net87619), .Z(net87627) );
  CNIVX3 U2970 ( .A(net87619), .Z(net87628) );
  CNIVX3 U2971 ( .A(net87619), .Z(net87629) );
  CNIVX3 U2972 ( .A(net87619), .Z(net87630) );
  CMX2XL U2973 ( .A0(\reg_mem[8][13] ), .A1(\reg_mem[9][13] ), .S(net87790), 
        .Z(n4296) );
  CMX2XL U2974 ( .A0(\reg_mem[0][5] ), .A1(\reg_mem[1][5] ), .S(net87790), .Z(
        n3954) );
  CMX2XL U2975 ( .A0(\reg_mem[2][5] ), .A1(\reg_mem[3][5] ), .S(net87790), .Z(
        n3953) );
  CMX2XL U2976 ( .A0(\reg_mem[0][17] ), .A1(\reg_mem[1][17] ), .S(net87795), 
        .Z(n4476) );
  CMX2XL U2977 ( .A0(\reg_mem[2][17] ), .A1(\reg_mem[3][17] ), .S(net87795), 
        .Z(n4475) );
  CMX2XL U2978 ( .A0(\reg_mem[16][16] ), .A1(\reg_mem[17][16] ), .S(net87790), 
        .Z(n4450) );
  CMX2XL U2979 ( .A0(\reg_mem[18][16] ), .A1(\reg_mem[19][16] ), .S(net87790), 
        .Z(n4449) );
  CMX2XL U2980 ( .A0(\reg_mem[20][16] ), .A1(\reg_mem[21][16] ), .S(net87790), 
        .Z(n4454) );
  CMX2XL U2981 ( .A0(\reg_mem[0][19] ), .A1(\reg_mem[1][19] ), .S(net87790), 
        .Z(n4564) );
  CMX2XL U2982 ( .A0(\reg_mem[0][20] ), .A1(\reg_mem[1][20] ), .S(net87790), 
        .Z(n4604) );
  CMX2XL U2983 ( .A0(\reg_mem[2][20] ), .A1(\reg_mem[3][20] ), .S(net87790), 
        .Z(n4603) );
  CMX2XL U2984 ( .A0(\reg_mem[0][7] ), .A1(\reg_mem[1][7] ), .S(net87790), .Z(
        n4042) );
  CMX2XL U2985 ( .A0(\reg_mem[0][10] ), .A1(\reg_mem[1][10] ), .S(net87790), 
        .Z(n4176) );
  CMX2XL U2986 ( .A0(\reg_mem[2][10] ), .A1(\reg_mem[3][10] ), .S(net87790), 
        .Z(n4175) );
  CMX2XL U2987 ( .A0(\reg_mem[8][10] ), .A1(\reg_mem[9][10] ), .S(net87790), 
        .Z(n4184) );
  CMX2XL U2988 ( .A0(\reg_mem[4][10] ), .A1(\reg_mem[5][10] ), .S(net87790), 
        .Z(n4180) );
  CMX2XL U2989 ( .A0(\reg_mem[12][10] ), .A1(\reg_mem[13][10] ), .S(net87790), 
        .Z(n4188) );
  CMX2XL U2990 ( .A0(\reg_mem[0][11] ), .A1(\reg_mem[1][11] ), .S(net87790), 
        .Z(net78097) );
  CMX2XL U2991 ( .A0(\reg_mem[16][10] ), .A1(\reg_mem[17][10] ), .S(net87790), 
        .Z(n4194) );
  CMX2XL U2992 ( .A0(\reg_mem[20][10] ), .A1(\reg_mem[21][10] ), .S(net87790), 
        .Z(n4198) );
  CMXI2X1 U2993 ( .A0(n2738), .A1(n2739), .S(n2169), .Z(n2743) );
  CMX2XL U2994 ( .A0(\reg_mem[20][7] ), .A1(\reg_mem[21][7] ), .S(net87790), 
        .Z(n4064) );
  CMXI2XL U2995 ( .A0(n4086), .A1(n4085), .S(net87803), .Z(n4088) );
  COND1X1 U2996 ( .A(n2454), .B(N30), .C(n2453), .Z(n2135) );
  CND2IX2 U2997 ( .B(n2067), .A(net87508), .Z(n3631) );
  CND2IXL U2998 ( .B(n3623), .A(n2568), .Z(n2577) );
  CND2X1 U2999 ( .A(n2067), .B(net87856), .Z(n3623) );
  CNIVX3 U3000 ( .A(n2076), .Z(n2105) );
  CND2X1 U3001 ( .A(N195), .B(n2140), .Z(n2666) );
  CIVXL U3002 ( .A(net87522), .Z(net87510) );
  CIVX2 U3003 ( .A(n1472), .Z(net87511) );
  CIVX1 U3004 ( .A(net83575), .Z(net87512) );
  CIVX1 U3005 ( .A(n1472), .Z(net87513) );
  CNIVX3 U3006 ( .A(net87513), .Z(net87524) );
  CNIVX2 U3007 ( .A(net87512), .Z(net87526) );
  COAN1X1 U3008 ( .A(n3641), .B(n3640), .C(n3639), .Z(n2065) );
  CND2X1 U3009 ( .A(n2065), .B(n3638), .Z(N299) );
  CND3XL U3010 ( .A(n3615), .B(n3614), .C(n3613), .Z(n3641) );
  CND2XL U3011 ( .A(n1533), .B(n3643), .Z(n3639) );
  CND2X1 U3012 ( .A(N199), .B(n2140), .Z(n3638) );
  CMXI2X1 U3013 ( .A0(n4138), .A1(n4137), .S(net87704), .Z(n4148) );
  CND2IX2 U3014 ( .B(n2448), .A(N32), .Z(n2452) );
  CIVX3 U3015 ( .A(n2038), .Z(n2180) );
  CMXI2XL U3016 ( .A0(n4008), .A1(n4007), .S(net87802), .Z(n4009) );
  CMXI2XL U3017 ( .A0(n4018), .A1(n4017), .S(net87803), .Z(n4019) );
  CMXI2XL U3018 ( .A0(n4000), .A1(n3999), .S(net87804), .Z(n4001) );
  CMXI2XL U3019 ( .A0(n3517), .A1(n3516), .S(n2089), .Z(n3519) );
  CMXI2XL U3020 ( .A0(\reg_mem[15][30] ), .A1(\reg_mem[31][30] ), .S(n2089), 
        .Z(n3599) );
  CMXI2XL U3021 ( .A0(\reg_mem[0][28] ), .A1(\reg_mem[16][28] ), .S(n2089), 
        .Z(n2554) );
  CMXI2XL U3022 ( .A0(n4669), .A1(n4699), .S(n2089), .Z(n2838) );
  CIVX2 U3023 ( .A(n2167), .Z(n2175) );
  CMXI2XL U3024 ( .A0(\reg_mem[11][29] ), .A1(\reg_mem[27][29] ), .S(n2086), 
        .Z(n2527) );
  CMXI2XL U3025 ( .A0(n4377), .A1(n4407), .S(n2098), .Z(n3045) );
  CND2IXL U3026 ( .B(n3653), .A(n3049), .Z(n3054) );
  CND2IXL U3027 ( .B(n3653), .A(n2837), .Z(n2842) );
  CMXI2X1 U3028 ( .A0(n2888), .A1(n1668), .S(n1480), .Z(n2896) );
  CMXI2XL U3029 ( .A0(n2911), .A1(n2910), .S(n2201), .Z(n2915) );
  CNR2X1 U3030 ( .A(n2825), .B(n2120), .Z(n2826) );
  CNR4X2 U3031 ( .A(n2821), .B(n2824), .C(n2823), .D(n2822), .Z(n2825) );
  CNIVX1 U3032 ( .A(net87239), .Z(net87275) );
  CMXI2XL U3033 ( .A0(n3125), .A1(n3124), .S(n2199), .Z(n3126) );
  CIVX2 U3034 ( .A(n2805), .Z(n2076) );
  CIVX1 U3035 ( .A(net79756), .Z(net87376) );
  CIVX1 U3036 ( .A(net79756), .Z(net87377) );
  CIVX1 U3037 ( .A(net79756), .Z(net87379) );
  CNIVX4 U3038 ( .A(n2053), .Z(n2069) );
  CNIVX1 U3039 ( .A(n2053), .Z(n2070) );
  CNIVX4 U3040 ( .A(net87374), .Z(net87385) );
  CNIVX4 U3041 ( .A(net87380), .Z(net87389) );
  CNIVX2 U3042 ( .A(net87378), .Z(net87392) );
  CNIVX4 U3043 ( .A(net87376), .Z(net87393) );
  CNIVX4 U3044 ( .A(net87376), .Z(net87394) );
  CNIVX4 U3045 ( .A(net87376), .Z(net87395) );
  CNIVX4 U3046 ( .A(net87377), .Z(net87397) );
  CNIVX4 U3047 ( .A(net87377), .Z(net87398) );
  CNIVX2 U3048 ( .A(net87377), .Z(net87399) );
  CNIVX2 U3049 ( .A(net87377), .Z(net87400) );
  CNIVX2 U3050 ( .A(net87378), .Z(net87402) );
  CNIVX3 U3051 ( .A(net87378), .Z(net87403) );
  CNIVX2 U3052 ( .A(net87379), .Z(net87405) );
  CNIVX4 U3053 ( .A(net87379), .Z(net87406) );
  CNIVX4 U3054 ( .A(net87379), .Z(net87407) );
  CMXI2XL U3055 ( .A0(\reg_mem[7][31] ), .A1(\reg_mem[23][31] ), .S(n2085), 
        .Z(n3646) );
  CMXI2XL U3056 ( .A0(\reg_mem[4][21] ), .A1(\reg_mem[20][21] ), .S(n2085), 
        .Z(n2859) );
  CMX2X1 U3057 ( .A0(\reg_mem[24][25] ), .A1(\reg_mem[8][25] ), .S(n1382), .Z(
        n2696) );
  CMXI2XL U3058 ( .A0(n2731), .A1(n2730), .S(n1532), .Z(n2747) );
  CIVX2 U3059 ( .A(net79770), .Z(net87234) );
  CMXI2X1 U3060 ( .A0(n2733), .A1(n2732), .S(n2187), .Z(n2737) );
  CMXI2XL U3061 ( .A0(\reg_mem[5][30] ), .A1(\reg_mem[21][30] ), .S(n2096), 
        .Z(n3627) );
  CMXI2XL U3062 ( .A0(\reg_mem[13][27] ), .A1(\reg_mem[29][27] ), .S(n2096), 
        .Z(n2591) );
  CMXI2XL U3063 ( .A0(n4664), .A1(n4694), .S(n2096), .Z(n2844) );
  CMXI2XL U3064 ( .A0(n4881), .A1(n4911), .S(n2096), .Z(n2674) );
  CMXI2X1 U3065 ( .A0(n3576), .A1(n1537), .S(n2198), .Z(n3577) );
  CMXI2XL U3066 ( .A0(n3617), .A1(n3616), .S(n2198), .Z(n3621) );
  CMXI2XL U3067 ( .A0(n3418), .A1(n3417), .S(n2198), .Z(n3422) );
  CMXI2XL U3068 ( .A0(n2879), .A1(n2878), .S(n2198), .Z(n2880) );
  CIVX1 U3069 ( .A(n2167), .Z(n2170) );
  CMXI2X1 U3070 ( .A0(n2735), .A1(n2734), .S(n1383), .Z(n2736) );
  CNIVX4 U3071 ( .A(regA[27]), .Z(n2071) );
  CIVX2 U3072 ( .A(net87251), .Z(net87231) );
  CIVX1 U3073 ( .A(net79770), .Z(net87235) );
  CIVXL U3074 ( .A(net79770), .Z(net87236) );
  CIVXL U3075 ( .A(net79770), .Z(net87237) );
  CIVXL U3076 ( .A(net79770), .Z(net87238) );
  CIVXL U3077 ( .A(net79770), .Z(net87239) );
  CNIVX4 U3078 ( .A(net87234), .Z(net87243) );
  CNIVX2 U3079 ( .A(net87241), .Z(net87251) );
  CNIVX2 U3080 ( .A(net87236), .Z(net87252) );
  CNIVX2 U3081 ( .A(net87236), .Z(net87253) );
  CNIVX2 U3082 ( .A(net87236), .Z(net87255) );
  CNIVX2 U3083 ( .A(net87236), .Z(net87256) );
  CNIVX2 U3084 ( .A(net87237), .Z(net87258) );
  CNIVX2 U3085 ( .A(net87237), .Z(net87260) );
  CNIVX2 U3086 ( .A(net87237), .Z(net87261) );
  CNIVX2 U3087 ( .A(net87238), .Z(net87263) );
  CNIVX2 U3088 ( .A(net87238), .Z(net87265) );
  CNIVX2 U3089 ( .A(net87238), .Z(net87266) );
  CNIVX2 U3090 ( .A(net87239), .Z(net87268) );
  CNIVX2 U3091 ( .A(net87239), .Z(net87269) );
  CNIVX2 U3092 ( .A(net87239), .Z(net87271) );
  CNIVX2 U3093 ( .A(net87237), .Z(net87272) );
  CNIVX2 U3094 ( .A(net87241), .Z(net87273) );
  CNIVX2 U3095 ( .A(net87241), .Z(net87276) );
  CIVXL U3096 ( .A(n2095), .Z(n2074) );
  CIVX2 U3097 ( .A(n2805), .Z(n2077) );
  CIVX2 U3098 ( .A(n2805), .Z(n2078) );
  CNIVX3 U3099 ( .A(n2077), .Z(n2085) );
  CNIVX4 U3100 ( .A(n2077), .Z(n2086) );
  CNIVX3 U3101 ( .A(n2076), .Z(n2087) );
  CNIVX3 U3102 ( .A(n2076), .Z(n2088) );
  CNIVX3 U3103 ( .A(n2078), .Z(n2089) );
  CNIVX4 U3104 ( .A(n2078), .Z(n2091) );
  CNIVX3 U3105 ( .A(n2079), .Z(n2092) );
  CNIVX3 U3106 ( .A(n2076), .Z(n2093) );
  CNIVX3 U3107 ( .A(n2079), .Z(n2095) );
  CNIVX3 U3108 ( .A(n2079), .Z(n2097) );
  CIVX2 U3109 ( .A(n1552), .Z(n2273) );
  CIVX2 U3110 ( .A(n2107), .Z(n2109) );
  CND2X1 U3111 ( .A(n2737), .B(net87233), .Z(n2111) );
  CND2X1 U3112 ( .A(n2736), .B(net87261), .Z(n2112) );
  CND2X1 U3113 ( .A(n2111), .B(n2112), .Z(n2113) );
  CNR2XL U3114 ( .A(n1533), .B(n2075), .Z(n2114) );
  CND2IXL U3115 ( .B(n3119), .A(n3118), .Z(alu_op_c[13]) );
  CANR1X2 U3116 ( .A(n2454), .B(n2452), .C(n2451), .Z(n2453) );
  CNIVX2 U3117 ( .A(n3695), .Z(n2115) );
  COR2XL U3118 ( .A(data_mem_rd_d), .B(i_type_wb), .Z(n2116) );
  COR2X1 U3119 ( .A(data_mem_rd_d), .B(i_type_wb), .Z(n2117) );
  CIVDX1 U3120 ( .A(n232), .Z0(net87043), .Z1(net87042) );
  CAN2XL U3121 ( .A(n1533), .B(n2828), .Z(n2120) );
  COND3XL U3122 ( .A(n2272), .B(n2789), .C(n2788), .D(n2787), .Z(n2828) );
  CND2X1 U3123 ( .A(n2815), .B(n1470), .Z(n2121) );
  CND2XL U3124 ( .A(n3748), .B(n3749), .Z(prog_count_c[7]) );
  CIVX1 U3125 ( .A(n2273), .Z(n2123) );
  CIVX1 U3126 ( .A(n2124), .Z(n2126) );
  CND2X1 U3127 ( .A(n219), .B(n204), .Z(n225) );
  CNR2IX2 U3128 ( .B(n3691), .A(N200), .Z(n3692) );
  CNR2X1 U3129 ( .A(n3686), .B(n2128), .Z(n3693) );
  CND2XL U3130 ( .A(n219), .B(n206), .Z(n226) );
  CND2X2 U3131 ( .A(n3562), .B(n3561), .Z(alu_op_c[1]) );
  CNR2X1 U3132 ( .A(net86999), .B(n2460), .Z(net80178) );
  CNR3X2 U3133 ( .A(n3685), .B(n3684), .C(n3683), .Z(n3686) );
  CANR2X1 U3134 ( .A(regc_addr_wb[3]), .B(n240), .C(regb_addr_wb[3]), .D(n2117), .Z(n208) );
  CIVXL U3135 ( .A(n2138), .Z(n3343) );
  CNR2XL U3136 ( .A(inst_fetch[3]), .B(inst_fetch[0]), .Z(n2460) );
  CAN2X1 U3137 ( .A(n1533), .B(n3687), .Z(n2128) );
  CND2XL U3138 ( .A(n3217), .B(n3216), .Z(alu_op_c[10]) );
  CND2IXL U3139 ( .B(net87385), .A(n2143), .Z(n2129) );
  CAN2X1 U3140 ( .A(net87275), .B(net87510), .Z(n2143) );
  CND2X1 U3141 ( .A(n2665), .B(n2666), .Z(N295) );
  CNIVXL U3142 ( .A(n239), .Z(n2210) );
  CNIVXL U3143 ( .A(n239), .Z(n2209) );
  CNIVXL U3144 ( .A(n239), .Z(n2212) );
  CNIVXL U3145 ( .A(n239), .Z(n2211) );
  CANR2XL U3146 ( .A(alu_op_c[2]), .B(n3750), .C(regA[2]), .D(n3739), .Z(n3528) );
  CAN2XL U3147 ( .A(n1533), .B(n3081), .Z(n2132) );
  CNR2XL U3148 ( .A(n3077), .B(n2132), .Z(n3078) );
  CND2XL U3149 ( .A(n3079), .B(n3078), .Z(N284) );
  CND2XL U3150 ( .A(n3007), .B(n3006), .Z(alu_op_c[16]) );
  CND2XL U3151 ( .A(n3148), .B(n3147), .Z(alu_op_c[12]) );
  CNR2X2 U3152 ( .A(n2147), .B(n3476), .Z(n2446) );
  CIVXL U3153 ( .A(n2167), .Z(n2133) );
  COND1XL U3154 ( .A(n2454), .B(N30), .C(n2042), .Z(n3329) );
  CND2XL U3155 ( .A(n2866), .B(n2867), .Z(N290) );
  CND2X1 U3156 ( .A(N192), .B(n3704), .Z(n2785) );
  CNR2IX1 U3157 ( .B(n5239), .A(n3332), .Z(n2147) );
  CNR2IX1 U3158 ( .B(N103), .A(n2123), .Z(n3287) );
  CND3X2 U3159 ( .A(n3699), .B(n3345), .C(n2153), .Z(n3563) );
  CANR2X1 U3160 ( .A(regc_addr_wb[0]), .B(n240), .C(regb_addr_wb[0]), .D(n241), 
        .Z(n229) );
  CANR2X1 U3161 ( .A(regc_addr_wb[4]), .B(n240), .C(regb_addr_wb[4]), .D(n2117), .Z(n207) );
  CND2XL U3162 ( .A(net87396), .B(n2083), .Z(n2796) );
  CNIVXL U3163 ( .A(net15031), .Z(net82869) );
  CNR2IX1 U3164 ( .B(n2136), .A(n2804), .Z(n2823) );
  CNR2XL U3165 ( .A(n2022), .B(n2069), .Z(n2136) );
  CNR2IXL U3166 ( .B(N104), .A(n2272), .Z(n3696) );
  CMXI2XL U3167 ( .A0(n2680), .A1(n2679), .S(n1469), .Z(n2684) );
  CND2XL U3168 ( .A(n2623), .B(n2622), .Z(n2629) );
  CNR3X1 U3169 ( .A(n229), .B(n230), .C(n5266), .Z(n196) );
  CNR3X1 U3170 ( .A(n231), .B(n230), .C(n5267), .Z(n194) );
  CANR2X1 U3171 ( .A(N170), .B(n3704), .C(N138), .D(n3701), .Z(n3559) );
  CND2IXL U3172 ( .B(n3474), .A(n3697), .Z(n3478) );
  CND2IXL U3173 ( .B(n3286), .A(N176), .Z(n3289) );
  CND2IXL U3174 ( .B(n3181), .A(N162), .Z(n2670) );
  CND2IXL U3175 ( .B(n3181), .A(N157), .Z(n2900) );
  CNR2IXL U3176 ( .B(n5238), .A(n3332), .Z(n3341) );
  CNR2IXL U3177 ( .B(N98), .A(n2272), .Z(n3520) );
  CNR2X1 U3178 ( .A(n3645), .B(n3644), .Z(n3687) );
  CNR2IXL U3179 ( .B(N114), .A(n2271), .Z(n2942) );
  CNR2IXL U3180 ( .B(N115), .A(n2115), .Z(n2907) );
  CND2XL U3181 ( .A(n2581), .B(n2580), .Z(n2587) );
  CND2IXL U3182 ( .B(n3694), .A(n2137), .Z(alu_op_c[31]) );
  CND2XL U3183 ( .A(N75), .B(n3697), .Z(n3183) );
  CND2XL U3184 ( .A(N78), .B(n3697), .Z(n3083) );
  CND3X1 U3185 ( .A(n2715), .B(n2714), .C(n2713), .Z(n2717) );
  CND2XL U3186 ( .A(N198), .B(n3704), .Z(n2544) );
  CANR1X1 U3187 ( .A(N167), .B(n3701), .C(n3635), .Z(n3637) );
  CMX2XL U3188 ( .A0(n1981), .A1(alu_op_c[18]), .S(n1533), .Z(N287) );
  CNR2IX1 U3189 ( .B(N120), .A(n2123), .Z(n2712) );
  CND2XL U3190 ( .A(n3528), .B(n3527), .Z(prog_count_c[2]) );
  CNR2IXL U3191 ( .B(n3526), .A(n3525), .Z(n3527) );
  CAN2XL U3192 ( .A(net87489), .B(inst_fetch[24]), .Z(net86659) );
  COND2XL U3193 ( .A(n2861), .B(n3681), .C(n2860), .D(n2129), .Z(n2862) );
  CMXI2XL U3194 ( .A0(\reg_mem[6][21] ), .A1(\reg_mem[22][21] ), .S(n2091), 
        .Z(n2858) );
  COND2XL U3195 ( .A(n3073), .B(n3681), .C(n3072), .D(n2129), .Z(n3074) );
  CMXI2XL U3196 ( .A0(\reg_mem[6][15] ), .A1(\reg_mem[22][15] ), .S(n2095), 
        .Z(n3070) );
  CNR2IXL U3197 ( .B(prog_count_ex[6]), .A(n3382), .Z(n2157) );
  COND4CXL U3198 ( .A(n5264), .B(n5238), .C(n5239), .D(opcode_ex[4]), .Z(n339)
         );
  CND2X1 U3199 ( .A(N168), .B(n3701), .Z(n3690) );
  CND2XL U3200 ( .A(opcode_ex[2]), .B(opcode_ex[5]), .Z(n2448) );
  CNR2IXL U3201 ( .B(prog_count_ex[4]), .A(n3430), .Z(n3383) );
  CANR2XL U3202 ( .A(alu_op_c[5]), .B(n3750), .C(regA[5]), .D(n3739), .Z(n3394) );
  CND2XL U3203 ( .A(N95), .B(n3697), .Z(n3688) );
  CND2XL U3204 ( .A(N127), .B(n2273), .Z(n3689) );
  CNR2X1 U3205 ( .A(opcode_ex[0]), .B(opcode_ex[4]), .Z(n2440) );
  CAN3X1 U3206 ( .A(prog_count_o[5]), .B(n3741), .C(n2154), .Z(n2155) );
  CNR2IXL U3207 ( .B(inst_fetch[29]), .A(net76768), .Z(n5233) );
  CNR2IXL U3208 ( .B(inst_fetch[30]), .A(net76768), .Z(n5234) );
  CNR2IXL U3209 ( .B(inst_fetch[31]), .A(net76768), .Z(n5236) );
  CND2IXL U3210 ( .B(n2069), .A(n2143), .Z(n3679) );
  CND2X1 U3211 ( .A(n1456), .B(n2143), .Z(n3649) );
  CAN2X1 U3212 ( .A(net87389), .B(n2142), .Z(n2139) );
  CANR1XL U3213 ( .A(N163), .B(n3701), .C(n2630), .Z(n2632) );
  CNIVX1 U3214 ( .A(net15031), .Z(net82859) );
  CNIVX1 U3215 ( .A(net15031), .Z(net82861) );
  CANR1XL U3216 ( .A(N164), .B(n3701), .C(n2621), .Z(n2623) );
  CND2X1 U3217 ( .A(n3633), .B(n3632), .Z(n3640) );
  CND2X1 U3218 ( .A(n2577), .B(n2576), .Z(n2584) );
  CND3XL U3219 ( .A(n3615), .B(n2561), .C(n2560), .Z(n2585) );
  CND2XL U3220 ( .A(n1533), .B(n2587), .Z(n2583) );
  CND2X1 U3221 ( .A(n228), .B(n204), .Z(n237) );
  CND2X1 U3222 ( .A(n228), .B(n200), .Z(n235) );
  CND2X1 U3223 ( .A(n228), .B(n192), .Z(n227) );
  CND2X1 U3224 ( .A(n2619), .B(n2618), .Z(n2626) );
  CND3XL U3225 ( .A(n3615), .B(n2603), .C(n2602), .Z(n2627) );
  CND2XL U3226 ( .A(n1533), .B(n2629), .Z(n2625) );
  CND3XL U3227 ( .A(n2843), .B(n2842), .C(n2841), .Z(n2864) );
  CANR1XL U3228 ( .A(n2139), .B(n2840), .C(n1533), .Z(n2841) );
  CND3XL U3229 ( .A(n3055), .B(n3054), .C(n3053), .Z(n3076) );
  CANR1XL U3230 ( .A(n2139), .B(n3052), .C(n1533), .Z(n3053) );
  CND3XL U3231 ( .A(n3067), .B(n3066), .C(n3065), .Z(n3075) );
  CNR2IX1 U3232 ( .B(n2813), .A(n2812), .Z(n2822) );
  CNR2IX1 U3233 ( .B(n2686), .A(n2646), .Z(n2662) );
  CNR2IXL U3234 ( .B(n1533), .A(n3694), .Z(n3691) );
  CND2XL U3235 ( .A(net87410), .B(net87533), .Z(n3604) );
  CND2IX1 U3236 ( .B(n2144), .A(n2826), .Z(N291) );
  CANR1XL U3237 ( .A(N74), .B(n3697), .C(n3215), .Z(n3216) );
  CND2X1 U3238 ( .A(n2909), .B(n2908), .Z(alu_op_c[19]) );
  CANR1XL U3239 ( .A(N83), .B(n3697), .C(n2907), .Z(n2908) );
  CANR1XL U3240 ( .A(N82), .B(n3697), .C(n2942), .Z(n2943) );
  CND2X1 U3241 ( .A(n3252), .B(n3251), .Z(alu_op_c[9]) );
  CANR1XL U3242 ( .A(N73), .B(n3697), .C(n3250), .Z(n3251) );
  CANR1XL U3243 ( .A(N80), .B(n3697), .C(n3005), .Z(n3006) );
  CANR1XL U3244 ( .A(N76), .B(n3697), .C(n3146), .Z(n3147) );
  CNR2IX1 U3245 ( .B(n3615), .A(n2899), .Z(n2904) );
  CND2X1 U3246 ( .A(N189), .B(n3704), .Z(n2905) );
  CNR2X1 U3247 ( .A(n207), .B(n208), .Z(n191) );
  CNR2X1 U3248 ( .A(n2502), .B(n2501), .Z(n2503) );
  CND3XL U3249 ( .A(n2498), .B(n2497), .C(n2496), .Z(n2502) );
  CNR3X1 U3250 ( .A(n229), .B(n230), .C(n231), .Z(n192) );
  CANR1XL U3251 ( .A(N173), .B(n3704), .C(n3433), .Z(n3434) );
  CANR1XL U3252 ( .A(N172), .B(n3704), .C(n1538), .Z(n3477) );
  CND2XL U3253 ( .A(N84), .B(n3697), .Z(n2901) );
  CND2XL U3254 ( .A(N89), .B(n3697), .Z(n2669) );
  CIVX2 U3255 ( .A(j_type_c), .Z(net76768) );
  CND2X1 U3256 ( .A(n3328), .B(n3327), .Z(alu_op_c[6]) );
  CANR1XL U3257 ( .A(N175), .B(n3704), .C(n3325), .Z(n3328) );
  CANR1XL U3258 ( .A(N70), .B(n3697), .C(n3326), .Z(n3327) );
  CANR1XL U3259 ( .A(N165), .B(n3701), .C(n2579), .Z(n2581) );
  CIVX2 U3260 ( .A(n3286), .Z(n3704) );
  CIVX1 U3261 ( .A(n2273), .Z(n2271) );
  CND2IX1 U3262 ( .B(n3345), .A(n2153), .Z(n3751) );
  CNR2IX1 U3263 ( .B(net76768), .A(n5242), .Z(n2145) );
  COND2XL U3264 ( .A(n2272), .B(n2974), .C(n3116), .D(n2973), .Z(n2976) );
  COND2XL U3265 ( .A(n2272), .B(n3117), .C(n3116), .D(n3115), .Z(n3119) );
  CND3XL U3266 ( .A(n2782), .B(n2781), .C(n2780), .Z(n2786) );
  CANR1XL U3267 ( .A(N66), .B(n3697), .C(n3522), .Z(n3523) );
  CNR2IX1 U3268 ( .B(n3521), .A(n3520), .Z(n3524) );
  CND3XL U3269 ( .A(n3690), .B(n3689), .C(n3688), .Z(n3694) );
  CND3XL U3270 ( .A(n3707), .B(n3706), .C(n3705), .Z(alu_op_c[8]) );
  CANR1XL U3271 ( .A(N177), .B(n3704), .C(n3703), .Z(n3705) );
  COND1XL U3272 ( .A(n5247), .B(net76768), .C(n5235), .Z(immi_val_c[15]) );
  CNR2IXL U3273 ( .B(N119), .A(n2272), .Z(n2779) );
  CND2X1 U3274 ( .A(n3689), .B(n3688), .Z(n3644) );
  CNIVX1 U3275 ( .A(n239), .Z(n2213) );
  CAN2XL U3276 ( .A(n3476), .B(n2153), .Z(n2146) );
  CNR2IXL U3277 ( .B(n2154), .A(n3563), .Z(n3393) );
  CNR2IX1 U3278 ( .B(n5217), .A(n2145), .Z(immi_val_c[0]) );
  CNR2IX1 U3279 ( .B(n5219), .A(n2145), .Z(immi_val_c[2]) );
  CNR2IX1 U3280 ( .B(n5220), .A(n2145), .Z(immi_val_c[3]) );
  CNR2IX1 U3281 ( .B(n5218), .A(n2145), .Z(immi_val_c[1]) );
  CNR2IX1 U3282 ( .B(n5221), .A(n2145), .Z(immi_val_c[4]) );
  CNR2IX1 U3283 ( .B(n5222), .A(n2145), .Z(immi_val_c[5]) );
  CNR2IX1 U3284 ( .B(n5223), .A(n2145), .Z(immi_val_c[6]) );
  CNR2IX1 U3285 ( .B(n5224), .A(n2145), .Z(immi_val_c[7]) );
  CNR2IX1 U3286 ( .B(n5225), .A(n2145), .Z(immi_val_c[8]) );
  CNR2IX1 U3287 ( .B(n5226), .A(n2145), .Z(immi_val_c[9]) );
  CNR2IX1 U3288 ( .B(n5227), .A(n2145), .Z(immi_val_c[10]) );
  CNR2X1 U3289 ( .A(n5251), .B(n2145), .Z(immi_val_c[11]) );
  CNR2X1 U3290 ( .A(n5250), .B(n2145), .Z(immi_val_c[12]) );
  CNR2X1 U3291 ( .A(n5249), .B(n2145), .Z(immi_val_c[13]) );
  CNR2X1 U3292 ( .A(n5248), .B(n2145), .Z(immi_val_c[14]) );
  CNIVX1 U3293 ( .A(n2203), .Z(n2208) );
  CNIVX1 U3294 ( .A(n2203), .Z(n2207) );
  CNIVX1 U3295 ( .A(n2203), .Z(n2206) );
  CNIVX1 U3296 ( .A(n2203), .Z(n2205) );
  CNIVX1 U3297 ( .A(n2203), .Z(n2204) );
  CANR1XL U3298 ( .A(N93), .B(n3697), .C(n2539), .Z(n2541) );
  CND2X1 U3299 ( .A(net87372), .B(n2142), .Z(n3667) );
  CND2IX1 U3300 ( .B(n3086), .A(n3085), .Z(alu_op_c[14]) );
  CND2IX1 U3301 ( .B(n3286), .A(N183), .Z(n3085) );
  CAN2XL U3302 ( .A(n1667), .B(net78793), .Z(net86675) );
  CND2XL U3303 ( .A(N184), .B(n2140), .Z(n3079) );
  CND2XL U3304 ( .A(N190), .B(n2140), .Z(n2867) );
  CNR2IXL U3305 ( .B(n3382), .A(n3699), .Z(n3386) );
  CNIVX1 U3306 ( .A(n242), .Z(n2274) );
  CNIVX1 U3307 ( .A(n242), .Z(n2275) );
  CNIVX1 U3308 ( .A(n242), .Z(n2277) );
  CNIVX1 U3309 ( .A(n242), .Z(n2276) );
  CNIVX1 U3310 ( .A(n242), .Z(n2278) );
  CND2X1 U3311 ( .A(inst_fetch[21]), .B(n5242), .Z(n5235) );
  CNR2IX1 U3312 ( .B(n3743), .A(n3742), .Z(n3744) );
  COND1XL U3313 ( .A(n3563), .B(prog_count_o[2]), .C(enable), .Z(n3481) );
  CENX1 U3314 ( .A(inst_fetch[30]), .B(regb_addr[3]), .Z(n2496) );
  CENX1 U3315 ( .A(inst_fetch[28]), .B(regb_addr[1]), .Z(n2497) );
  CMX2X1 U3316 ( .A0(\reg_mem[0][0] ), .A1(\reg_mem[1][0] ), .S(net87799), .Z(
        n3758) );
  CMX2X1 U3317 ( .A0(\reg_mem[0][3] ), .A1(\reg_mem[1][3] ), .S(net87804), .Z(
        n3878) );
  CMX2X1 U3318 ( .A0(\reg_mem[0][14] ), .A1(\reg_mem[1][14] ), .S(net87790), 
        .Z(n4328) );
  CMX2X1 U3319 ( .A0(\reg_mem[0][23] ), .A1(\reg_mem[1][23] ), .S(net87797), 
        .Z(n4772) );
  CMX2X1 U3320 ( .A0(\reg_mem[16][1] ), .A1(\reg_mem[17][1] ), .S(net87800), 
        .Z(n3820) );
  CMX2X1 U3321 ( .A0(\reg_mem[16][5] ), .A1(\reg_mem[17][5] ), .S(net87795), 
        .Z(n3972) );
  CMX2X1 U3322 ( .A0(\reg_mem[16][8] ), .A1(\reg_mem[17][8] ), .S(net87790), 
        .Z(n4106) );
  CMX2X1 U3323 ( .A0(\reg_mem[16][12] ), .A1(\reg_mem[17][12] ), .S(net87790), 
        .Z(n4270) );
  CMX2X1 U3324 ( .A0(\reg_mem[4][1] ), .A1(\reg_mem[5][1] ), .S(net87798), .Z(
        n3806) );
  CMX2X1 U3325 ( .A0(\reg_mem[4][2] ), .A1(\reg_mem[5][2] ), .S(net87802), .Z(
        n3850) );
  CMX2X1 U3326 ( .A0(\reg_mem[4][3] ), .A1(\reg_mem[5][3] ), .S(net87804), .Z(
        n3882) );
  CMX2X1 U3327 ( .A0(\reg_mem[4][4] ), .A1(\reg_mem[5][4] ), .S(net87797), .Z(
        n3926) );
  CMX2X1 U3328 ( .A0(\reg_mem[4][7] ), .A1(\reg_mem[5][7] ), .S(net87802), .Z(
        n4046) );
  CMX2X1 U3329 ( .A0(\reg_mem[4][9] ), .A1(\reg_mem[5][9] ), .S(net87790), .Z(
        n4136) );
  CMX2X1 U3330 ( .A0(\reg_mem[4][14] ), .A1(\reg_mem[5][14] ), .S(net87804), 
        .Z(n4332) );
  CMX2X1 U3331 ( .A0(\reg_mem[4][16] ), .A1(\reg_mem[5][16] ), .S(net87795), 
        .Z(n4436) );
  CMX2X1 U3332 ( .A0(\reg_mem[4][23] ), .A1(\reg_mem[5][23] ), .S(net87809), 
        .Z(n4776) );
  CMX2X1 U3333 ( .A0(\reg_mem[20][1] ), .A1(\reg_mem[21][1] ), .S(net87799), 
        .Z(n3824) );
  CMX2X1 U3334 ( .A0(\reg_mem[20][8] ), .A1(\reg_mem[21][8] ), .S(net87798), 
        .Z(n4110) );
  CMX2X1 U3335 ( .A0(\reg_mem[20][11] ), .A1(\reg_mem[21][11] ), .S(net87799), 
        .Z(n4232) );
  CMX2X1 U3336 ( .A0(\reg_mem[20][17] ), .A1(\reg_mem[21][17] ), .S(net87803), 
        .Z(n4498) );
  CMX2X1 U3337 ( .A0(\reg_mem[8][0] ), .A1(\reg_mem[9][0] ), .S(net87790), .Z(
        n3766) );
  CMX2X1 U3338 ( .A0(\reg_mem[8][4] ), .A1(\reg_mem[9][4] ), .S(net87803), .Z(
        n3930) );
  CMX2X1 U3339 ( .A0(\reg_mem[8][16] ), .A1(\reg_mem[9][16] ), .S(net87790), 
        .Z(n4440) );
  CMX2X1 U3340 ( .A0(\reg_mem[8][17] ), .A1(\reg_mem[9][17] ), .S(net87791), 
        .Z(n4484) );
  CMX2X1 U3341 ( .A0(\reg_mem[12][0] ), .A1(\reg_mem[13][0] ), .S(net87802), 
        .Z(n3770) );
  CMX2X1 U3342 ( .A0(\reg_mem[12][1] ), .A1(\reg_mem[13][1] ), .S(net87802), 
        .Z(n3814) );
  CMX2X1 U3343 ( .A0(\reg_mem[12][3] ), .A1(\reg_mem[13][3] ), .S(net87794), 
        .Z(n3890) );
  CMX2X1 U3344 ( .A0(\reg_mem[12][4] ), .A1(\reg_mem[13][4] ), .S(net87806), 
        .Z(n3934) );
  CMX2X1 U3345 ( .A0(\reg_mem[12][7] ), .A1(\reg_mem[13][7] ), .S(net87797), 
        .Z(n4054) );
  CMX2X1 U3346 ( .A0(\reg_mem[12][8] ), .A1(\reg_mem[13][8] ), .S(net87803), 
        .Z(n4100) );
  CMX2X1 U3347 ( .A0(\reg_mem[12][16] ), .A1(\reg_mem[13][16] ), .S(net87804), 
        .Z(n4444) );
  CMX2X1 U3348 ( .A0(\reg_mem[12][17] ), .A1(\reg_mem[13][17] ), .S(net87809), 
        .Z(n4488) );
  CMX2X1 U3349 ( .A0(\reg_mem[12][18] ), .A1(\reg_mem[13][18] ), .S(net87795), 
        .Z(n4532) );
  CMX2X1 U3350 ( .A0(\reg_mem[12][19] ), .A1(\reg_mem[13][19] ), .S(net87795), 
        .Z(n4574) );
  CMX2X1 U3351 ( .A0(\reg_mem[0][29] ), .A1(\reg_mem[1][29] ), .S(net87797), 
        .Z(n5068) );
  CMX2X1 U3352 ( .A0(\reg_mem[16][23] ), .A1(\reg_mem[17][23] ), .S(net87798), 
        .Z(n4790) );
  CMX2X1 U3353 ( .A0(\reg_mem[16][28] ), .A1(\reg_mem[17][28] ), .S(net87795), 
        .Z(n5040) );
  CMX2X1 U3354 ( .A0(\reg_mem[16][29] ), .A1(\reg_mem[17][29] ), .S(net87794), 
        .Z(n5088) );
  CMX2X1 U3355 ( .A0(\reg_mem[16][30] ), .A1(\reg_mem[17][30] ), .S(net87806), 
        .Z(n5134) );
  CMX2X1 U3356 ( .A0(\reg_mem[4][28] ), .A1(\reg_mem[5][28] ), .S(net87803), 
        .Z(n5026) );
  CMX2X1 U3357 ( .A0(\reg_mem[12][30] ), .A1(\reg_mem[13][30] ), .S(net87809), 
        .Z(n5128) );
  CMX2X1 U3358 ( .A0(\reg_mem[20][23] ), .A1(\reg_mem[21][23] ), .S(net87809), 
        .Z(n4794) );
  CMX2X1 U3359 ( .A0(\reg_mem[20][28] ), .A1(\reg_mem[21][28] ), .S(net87807), 
        .Z(n5044) );
  CMX2X1 U3360 ( .A0(\reg_mem[20][30] ), .A1(\reg_mem[21][30] ), .S(net87806), 
        .Z(n5138) );
  CMX2X1 U3361 ( .A0(\reg_mem[8][23] ), .A1(\reg_mem[9][23] ), .S(net87807), 
        .Z(n4780) );
  CMX2X1 U3362 ( .A0(\reg_mem[0][30] ), .A1(\reg_mem[1][30] ), .S(net87798), 
        .Z(n5116) );
  CMX2X1 U3363 ( .A0(\reg_mem[12][23] ), .A1(\reg_mem[13][23] ), .S(net87794), 
        .Z(n4784) );
  CMX2X1 U3364 ( .A0(\reg_mem[12][29] ), .A1(\reg_mem[13][29] ), .S(net87798), 
        .Z(n5080) );
  CMX2X1 U3365 ( .A0(\reg_mem[4][30] ), .A1(\reg_mem[5][30] ), .S(net87793), 
        .Z(n5120) );
  CMXI2X1 U3366 ( .A0(n2508), .A1(n2507), .S(n2180), .Z(n2512) );
  CMX2X1 U3367 ( .A0(\reg_mem[2][0] ), .A1(\reg_mem[3][0] ), .S(net87799), .Z(
        n3757) );
  CMX2X1 U3368 ( .A0(\reg_mem[2][1] ), .A1(\reg_mem[3][1] ), .S(net87802), .Z(
        n3801) );
  CMX2X1 U3369 ( .A0(\reg_mem[2][4] ), .A1(\reg_mem[3][4] ), .S(net87804), .Z(
        n3921) );
  CMX2X1 U3370 ( .A0(\reg_mem[2][9] ), .A1(\reg_mem[3][9] ), .S(net87790), .Z(
        n4131) );
  CMX2X1 U3371 ( .A0(\reg_mem[2][19] ), .A1(\reg_mem[3][19] ), .S(net87793), 
        .Z(n4563) );
  CMX2X1 U3372 ( .A0(\reg_mem[2][23] ), .A1(\reg_mem[3][23] ), .S(net87807), 
        .Z(n4771) );
  CMX2X1 U3373 ( .A0(\reg_mem[18][1] ), .A1(\reg_mem[19][1] ), .S(net87799), 
        .Z(n3819) );
  CMX2X1 U3374 ( .A0(\reg_mem[18][6] ), .A1(\reg_mem[19][6] ), .S(net87797), 
        .Z(n4015) );
  CMX2X1 U3375 ( .A0(\reg_mem[18][9] ), .A1(\reg_mem[19][9] ), .S(net87790), 
        .Z(n4149) );
  CMX2X1 U3376 ( .A0(\reg_mem[18][12] ), .A1(\reg_mem[19][12] ), .S(net87790), 
        .Z(n4269) );
  CMX2X1 U3377 ( .A0(\reg_mem[18][20] ), .A1(\reg_mem[19][20] ), .S(net87809), 
        .Z(n4621) );
  CMX2X1 U3378 ( .A0(\reg_mem[10][1] ), .A1(\reg_mem[11][1] ), .S(net87797), 
        .Z(n3809) );
  CMX2X1 U3379 ( .A0(\reg_mem[10][3] ), .A1(\reg_mem[11][3] ), .S(net87804), 
        .Z(n3885) );
  CMX2X1 U3380 ( .A0(\reg_mem[10][5] ), .A1(\reg_mem[11][5] ), .S(net87803), 
        .Z(n3961) );
  CMX2X1 U3381 ( .A0(\reg_mem[10][14] ), .A1(\reg_mem[11][14] ), .S(net87795), 
        .Z(n4335) );
  CMX2X1 U3382 ( .A0(\reg_mem[10][16] ), .A1(\reg_mem[11][16] ), .S(net87800), 
        .Z(n4439) );
  CMX2X1 U3383 ( .A0(\reg_mem[10][17] ), .A1(\reg_mem[11][17] ), .S(net87795), 
        .Z(n4483) );
  CMX2X1 U3384 ( .A0(\reg_mem[10][20] ), .A1(\reg_mem[11][20] ), .S(net87795), 
        .Z(n4611) );
  CMX2X1 U3385 ( .A0(\reg_mem[2][27] ), .A1(\reg_mem[3][27] ), .S(net87790), 
        .Z(n4983) );
  CMX2X1 U3386 ( .A0(\reg_mem[10][30] ), .A1(\reg_mem[11][30] ), .S(net87793), 
        .Z(n5123) );
  CMX2X1 U3387 ( .A0(\reg_mem[18][23] ), .A1(\reg_mem[19][23] ), .S(net87804), 
        .Z(n4789) );
  CMX2X1 U3388 ( .A0(\reg_mem[18][28] ), .A1(\reg_mem[19][28] ), .S(net87802), 
        .Z(n5039) );
  CMX2X1 U3389 ( .A0(\reg_mem[10][23] ), .A1(\reg_mem[11][23] ), .S(net87809), 
        .Z(n4779) );
  CMX2X1 U3390 ( .A0(\reg_mem[10][24] ), .A1(\reg_mem[11][24] ), .S(net87790), 
        .Z(n4823) );
  CMX2X1 U3391 ( .A0(\reg_mem[2][30] ), .A1(\reg_mem[3][30] ), .S(net87791), 
        .Z(n5115) );
  CMX2X1 U3392 ( .A0(\reg_mem[10][31] ), .A1(\reg_mem[11][31] ), .S(net87790), 
        .Z(n5173) );
  CENX1 U3393 ( .A(inst_fetch[29]), .B(regb_addr[2]), .Z(n2498) );
  COND1XL U3394 ( .A(n2154), .B(n3563), .C(enable), .Z(n3392) );
  CND4X1 U3395 ( .A(n3342), .B(n3341), .C(n3340), .D(n3339), .Z(n3345) );
  CNR2X1 U3396 ( .A(n3334), .B(n3333), .Z(n3340) );
  CNR2X1 U3397 ( .A(n3338), .B(n3337), .Z(n3339) );
  CANR1XL U3398 ( .A(n2493), .B(n2492), .C(inst_fetch[27]), .Z(n2494) );
  CNR2X1 U3399 ( .A(regb_addr[3]), .B(regb_addr[4]), .Z(n2492) );
  CNR2X1 U3400 ( .A(regb_addr[1]), .B(regb_addr[2]), .Z(n2493) );
  CEOXL U3401 ( .A(n2157), .B(prog_count_ex[7]), .Z(n3285) );
  CND3XL U3402 ( .A(n2459), .B(n2458), .C(n2457), .Z(alu_op_c[0]) );
  CANR2XL U3403 ( .A(n3704), .B(N169), .C(N137), .D(n3701), .Z(n2459) );
  CND2XL U3404 ( .A(N96), .B(n2273), .Z(n2458) );
  CANR2XL U3405 ( .A(N128), .B(n3476), .C(N64), .D(n3697), .Z(n2457) );
  COR2XL U3406 ( .A(i_type_wb), .B(n240), .Z(n2203) );
  CMX2GXL U3407 ( .GN(n3563), .A0(prog_count_o[4]), .A1(n3438), .S(
        prog_count_o[3]), .Z(n3439) );
  CNR2X1 U3408 ( .A(n3480), .B(prog_count_o[4]), .Z(n3438) );
  CNR2XL U3409 ( .A(n2272), .B(n2538), .Z(n2539) );
  CNR2XL U3410 ( .A(n2271), .B(n2578), .Z(n2579) );
  CNR2IXL U3411 ( .B(n2109), .A(n3751), .Z(n3564) );
  CNR2IXL U3412 ( .B(n1388), .A(n3751), .Z(n3752) );
  CNR2XL U3413 ( .A(prog_count_ex[2]), .B(n3699), .Z(n3522) );
  CNR2IXL U3414 ( .B(N129), .A(n3699), .Z(n3560) );
  CNR2IXL U3415 ( .B(regA[4]), .A(n3751), .Z(n3440) );
  CAN3X2 U3416 ( .A(prog_count_o[2]), .B(prog_count_o[3]), .C(prog_count_o[4]), 
        .Z(n2154) );
  CNR2XL U3417 ( .A(prog_count_ex[5]), .B(n3383), .Z(n3384) );
  CNR2X1 U3418 ( .A(opcode_ext_ex[5]), .B(opcode_ext_ex[6]), .Z(n3336) );
  CNR2X1 U3419 ( .A(opcode_ext_ex[8]), .B(opcode_ext_ex[9]), .Z(n3335) );
  CND3XL U3420 ( .A(n3396), .B(n3395), .C(n3394), .Z(prog_count_c[5]) );
  CND2XL U3421 ( .A(prog_count_ex[5]), .B(n3383), .Z(n3382) );
  CANR3XL U3422 ( .A(n341), .B(n342), .C(opcode_ex[4]), .D(opcode_ex[0]), .Z(
        n340) );
  CND3XL U3423 ( .A(opcode_ex[1]), .B(opcode_ex[5]), .C(opcode_ex[2]), .Z(n341) );
  CND3XL U3424 ( .A(n5264), .B(n5240), .C(n5246), .Z(n342) );
  CND2XL U3425 ( .A(enable), .B(n3563), .Z(n3753) );
  CND2XL U3426 ( .A(prog_count_ex[2]), .B(prog_count_ex[3]), .Z(n3430) );
  CND3XL U3427 ( .A(n3348), .B(n3347), .C(n3346), .Z(prog_count_c[6]) );
  CND3XL U3428 ( .A(n3756), .B(n3755), .C(n3754), .Z(prog_count_c[0]) );
  CANR1XL U3429 ( .A(N22), .B(n3753), .C(n3752), .Z(n3754) );
  CND2XL U3430 ( .A(alu_op_c[0]), .B(n3750), .Z(n3756) );
  CND3XL U3431 ( .A(n3567), .B(n3566), .C(n3565), .Z(prog_count_c[1]) );
  CANR1XL U3432 ( .A(N23), .B(n3753), .C(n3564), .Z(n3565) );
  CND2XL U3433 ( .A(alu_op_c[1]), .B(n3750), .Z(n3567) );
  CND2XL U3434 ( .A(enable), .B(n3344), .Z(n3437) );
  CND3XL U3435 ( .A(n3443), .B(n3442), .C(n3441), .Z(prog_count_c[4]) );
  CANR3XL U3436 ( .A(prog_count_o[4]), .B(n3481), .C(n3440), .D(n3439), .Z(
        n3441) );
  CND2X1 U3437 ( .A(net86675), .B(n5215), .Z(n5216) );
  CNR2IX1 U3438 ( .B(inst_fetch[24]), .A(net76768), .Z(n5228) );
  CNR2IX1 U3439 ( .B(inst_fetch[25]), .A(net76768), .Z(n5229) );
  CNR2IX1 U3440 ( .B(inst_fetch[26]), .A(net76768), .Z(n5230) );
  CNR2IXL U3441 ( .B(inst_fetch[27]), .A(net76768), .Z(n5231) );
  CNR2IX1 U3442 ( .B(inst_fetch[28]), .A(net76768), .Z(n5232) );
  CND2X1 U3443 ( .A(n2500), .B(n2499), .Z(n2501) );
  CENX1 U3444 ( .A(inst_fetch[31]), .B(regb_addr[4]), .Z(n2499) );
  CND4XL U3445 ( .A(opcode_ex[4]), .B(opcode_ex[0]), .C(n2156), .D(n5239), .Z(
        n2500) );
  CND2X1 U3446 ( .A(opcode_ext_ex[4]), .B(opcode_ext_ex[3]), .Z(n3333) );
  CND2X1 U3447 ( .A(opcode_ext_ex[2]), .B(opcode_ext_ex[0]), .Z(n3334) );
  CEOXL U3448 ( .A(prog_count_ex[2]), .B(prog_count_ex[3]), .Z(n3475) );
  CNR2IX1 U3449 ( .B(n3747), .A(n3746), .Z(n3748) );
  CND2X1 U3450 ( .A(n3487), .B(n3486), .Z(prog_count_c[3]) );
  CNR2IX1 U3451 ( .B(n3485), .A(n3484), .Z(n3486) );
  CNR2IXL U3452 ( .B(prog_count_ex[7]), .A(n3699), .Z(n3700) );
  CND4X1 U3453 ( .A(n98), .B(n100), .C(opcode_mem[0]), .D(n249), .Z(n242) );
  CNR2X1 U3454 ( .A(n99), .B(n5268), .Z(n249) );
  CNR2X1 U3455 ( .A(opcode_mem[1]), .B(opcode_mem[0]), .Z(n248) );
  CNR2IX1 U3456 ( .B(opcode_mem[1]), .A(n2274), .Z(data_mem_rd_o) );
  CNR2X1 U3457 ( .A(opcode_mem[1]), .B(n2274), .Z(data_mem_wr_o) );
  CNR2IX1 U3458 ( .B(regB_mem[0]), .A(n2276), .Z(data_mem_wdata_o[0]) );
  CNR2IX1 U3459 ( .B(regB_mem[1]), .A(n2275), .Z(data_mem_wdata_o[1]) );
  CNR2IX1 U3460 ( .B(regB_mem[2]), .A(n2274), .Z(data_mem_wdata_o[2]) );
  CNR2IX1 U3461 ( .B(regB_mem[3]), .A(n2274), .Z(data_mem_wdata_o[3]) );
  CNR2IX1 U3462 ( .B(regB_mem[4]), .A(n2274), .Z(data_mem_wdata_o[4]) );
  CNR2IX1 U3463 ( .B(regB_mem[5]), .A(n2274), .Z(data_mem_wdata_o[5]) );
  CNR2IX1 U3464 ( .B(regB_mem[6]), .A(n2274), .Z(data_mem_wdata_o[6]) );
  CNR2IX1 U3465 ( .B(regB_mem[7]), .A(n2274), .Z(data_mem_wdata_o[7]) );
  CNR2IX1 U3466 ( .B(regB_mem[8]), .A(n2274), .Z(data_mem_wdata_o[8]) );
  CNR2IX1 U3467 ( .B(regB_mem[9]), .A(n2274), .Z(data_mem_wdata_o[9]) );
  CNR2IX1 U3468 ( .B(regB_mem[10]), .A(n2276), .Z(data_mem_wdata_o[10]) );
  CNR2IX1 U3469 ( .B(regB_mem[11]), .A(n2276), .Z(data_mem_wdata_o[11]) );
  CNR2IX1 U3470 ( .B(regB_mem[12]), .A(n2276), .Z(data_mem_wdata_o[12]) );
  CNR2IX1 U3471 ( .B(regB_mem[13]), .A(n2276), .Z(data_mem_wdata_o[13]) );
  CNR2IX1 U3472 ( .B(regB_mem[14]), .A(n2276), .Z(data_mem_wdata_o[14]) );
  CNR2IX1 U3473 ( .B(regB_mem[15]), .A(n2275), .Z(data_mem_wdata_o[15]) );
  CNR2IX1 U3474 ( .B(regB_mem[16]), .A(n2275), .Z(data_mem_wdata_o[16]) );
  CNR2IX1 U3475 ( .B(regB_mem[17]), .A(n2275), .Z(data_mem_wdata_o[17]) );
  CNR2IX1 U3476 ( .B(regB_mem[18]), .A(n2275), .Z(data_mem_wdata_o[18]) );
  CNR2IX1 U3477 ( .B(regB_mem[19]), .A(n2275), .Z(data_mem_wdata_o[19]) );
  CNR2IX1 U3478 ( .B(regB_mem[20]), .A(n2275), .Z(data_mem_wdata_o[20]) );
  CNR2IX1 U3479 ( .B(regB_mem[21]), .A(n2275), .Z(data_mem_wdata_o[21]) );
  CNR2IX1 U3480 ( .B(regB_mem[22]), .A(n2275), .Z(data_mem_wdata_o[22]) );
  CNR2IX1 U3481 ( .B(regB_mem[23]), .A(n2275), .Z(data_mem_wdata_o[23]) );
  CNR2IX1 U3482 ( .B(regB_mem[24]), .A(n2275), .Z(data_mem_wdata_o[24]) );
  CNR2IX1 U3483 ( .B(regB_mem[25]), .A(n2275), .Z(data_mem_wdata_o[25]) );
  CNR2IX1 U3484 ( .B(regB_mem[26]), .A(n2275), .Z(data_mem_wdata_o[26]) );
  CNR2IX1 U3485 ( .B(regB_mem[27]), .A(n2275), .Z(data_mem_wdata_o[27]) );
  CNR2IX1 U3486 ( .B(regB_mem[28]), .A(n2274), .Z(data_mem_wdata_o[28]) );
  CNR2IX1 U3487 ( .B(regB_mem[29]), .A(n2274), .Z(data_mem_wdata_o[29]) );
  CNR2IX1 U3488 ( .B(regB_mem[30]), .A(n2274), .Z(data_mem_wdata_o[30]) );
  CNR2IX1 U3489 ( .B(regB_mem[31]), .A(n2274), .Z(data_mem_wdata_o[31]) );
  CNR2IX1 U3490 ( .B(alu_op[0]), .A(n2278), .Z(data_mem_addr_o[0]) );
  CNR2IX1 U3491 ( .B(alu_op[1]), .A(n2277), .Z(data_mem_addr_o[1]) );
  CNR2IX1 U3492 ( .B(alu_op[2]), .A(n2277), .Z(data_mem_addr_o[2]) );
  CNR2IX1 U3493 ( .B(alu_op[3]), .A(n2276), .Z(data_mem_addr_o[3]) );
  CNR2IX1 U3494 ( .B(alu_op[4]), .A(n2276), .Z(data_mem_addr_o[4]) );
  CNR2IX1 U3495 ( .B(alu_op[5]), .A(n2276), .Z(data_mem_addr_o[5]) );
  CNR2IX1 U3496 ( .B(alu_op[6]), .A(n2276), .Z(data_mem_addr_o[6]) );
  CNR2IX1 U3497 ( .B(alu_op[7]), .A(n2276), .Z(data_mem_addr_o[7]) );
  CNR2IX1 U3498 ( .B(alu_op[8]), .A(n2276), .Z(data_mem_addr_o[8]) );
  CNR2IX1 U3499 ( .B(alu_op[9]), .A(n2276), .Z(data_mem_addr_o[9]) );
  CNR2IX1 U3500 ( .B(alu_op[10]), .A(n2278), .Z(data_mem_addr_o[10]) );
  CNR2IX1 U3501 ( .B(alu_op[11]), .A(n2278), .Z(data_mem_addr_o[11]) );
  CNR2IX1 U3502 ( .B(alu_op[12]), .A(n2278), .Z(data_mem_addr_o[12]) );
  CNR2IX1 U3503 ( .B(alu_op[13]), .A(n2278), .Z(data_mem_addr_o[13]) );
  CNR2IX1 U3504 ( .B(alu_op[14]), .A(n2278), .Z(data_mem_addr_o[14]) );
  CNR2IX1 U3505 ( .B(alu_op[15]), .A(n2278), .Z(data_mem_addr_o[15]) );
  CNR2IX1 U3506 ( .B(alu_op[16]), .A(n2278), .Z(data_mem_addr_o[16]) );
  CNR2IX1 U3507 ( .B(alu_op[17]), .A(n2278), .Z(data_mem_addr_o[17]) );
  CNR2IX1 U3508 ( .B(alu_op[18]), .A(n2278), .Z(data_mem_addr_o[18]) );
  CNR2IX1 U3509 ( .B(alu_op[19]), .A(n2277), .Z(data_mem_addr_o[19]) );
  CNR2IX1 U3510 ( .B(alu_op[20]), .A(n2277), .Z(data_mem_addr_o[20]) );
  CNR2IX1 U3511 ( .B(alu_op[21]), .A(n2277), .Z(data_mem_addr_o[21]) );
  CNR2IX1 U3512 ( .B(alu_op[22]), .A(n2277), .Z(data_mem_addr_o[22]) );
  CNR2IX1 U3513 ( .B(alu_op[23]), .A(n2277), .Z(data_mem_addr_o[23]) );
  CNR2IX1 U3514 ( .B(alu_op[24]), .A(n2277), .Z(data_mem_addr_o[24]) );
  CNR2IX1 U3515 ( .B(alu_op[25]), .A(n2277), .Z(data_mem_addr_o[25]) );
  CNR2IX1 U3516 ( .B(alu_op[26]), .A(n2277), .Z(data_mem_addr_o[26]) );
  CNR2IX1 U3517 ( .B(alu_op[27]), .A(n2277), .Z(data_mem_addr_o[27]) );
  CNR2IX1 U3518 ( .B(alu_op[28]), .A(n2277), .Z(data_mem_addr_o[28]) );
  CNR2IX1 U3519 ( .B(alu_op[29]), .A(n2277), .Z(data_mem_addr_o[29]) );
  CNR2IX1 U3520 ( .B(alu_op[30]), .A(n2277), .Z(data_mem_addr_o[30]) );
  CNR2IX1 U3521 ( .B(alu_op[31]), .A(n2276), .Z(data_mem_addr_o[31]) );
  CND2IXL U3522 ( .B(n3286), .A(N193), .Z(n2716) );
  CND2IXL U3523 ( .B(\dp_cluster_0/N57 ), .A(n2146), .Z(n3348) );
  CND2IXL U3524 ( .B(\dp_cluster_0/N62 ), .A(n2146), .Z(n3566) );
  CND2IXL U3525 ( .B(n1541), .A(n2146), .Z(n3755) );
  CND2IXL U3526 ( .B(n3286), .A(N180), .Z(n3185) );
  CND2XL U3527 ( .A(N196), .B(n3704), .Z(n2628) );
  CND2X1 U3528 ( .A(N197), .B(n2140), .Z(n2582) );
  CIVX2 U3529 ( .A(n2173), .Z(n2162) );
  CND2IXL U3530 ( .B(n1555), .A(n2146), .Z(n3747) );
  CIVXL U3531 ( .A(net88101), .Z(net76653) );
  CND2IXL U3532 ( .B(n1409), .A(n2146), .Z(n3526) );
  CND2IXL U3533 ( .B(n1556), .A(n2146), .Z(n3396) );
  CANR1X1 U3534 ( .A(inst_fetch[3]), .B(net78797), .C(inst_fetch[2]), .Z(n2163) );
  CIVX2 U3535 ( .A(n2169), .Z(n2166) );
  CNR2IX1 U3536 ( .B(n3693), .A(n3692), .Z(N300) );
  CNR2IX1 U3537 ( .B(n2694), .A(n2693), .Z(n2704) );
  CMXI2XL U3538 ( .A0(n2638), .A1(n2637), .S(net87272), .Z(n2639) );
  COND3X1 U3539 ( .A(n2585), .B(n2584), .C(n2582), .D(n2583), .Z(N297) );
  CNR4X2 U3540 ( .A(n2663), .B(n2660), .C(n2661), .D(n2662), .Z(n2664) );
  CND2X2 U3541 ( .A(net87488), .B(inst_fetch[27]), .Z(net79756) );
  CMXI2XL U3542 ( .A0(n3379), .A1(n3380), .S(n3615), .Z(N275) );
  CMXI2XL U3543 ( .A0(n3518), .A1(n3519), .S(n3615), .Z(N272) );
  CMXI2XL U3544 ( .A0(n3427), .A1(n3428), .S(n3615), .Z(N274) );
  CMXI2XL U3545 ( .A0(n3248), .A1(n3249), .S(n3615), .Z(N279) );
  CND2X2 U3546 ( .A(n2504), .B(n2503), .Z(n3615) );
  CIVX2 U3547 ( .A(n2167), .Z(n2171) );
  CIVX2 U3548 ( .A(n2167), .Z(n2173) );
  CIVX2 U3549 ( .A(n2167), .Z(n2174) );
  CIVX2 U3550 ( .A(n2175), .Z(n2176) );
  CIVX2 U3551 ( .A(n2038), .Z(n2177) );
  CIVX2 U3552 ( .A(n2168), .Z(n2178) );
  CIVX2 U3553 ( .A(n2038), .Z(n2179) );
  CIVX2 U3554 ( .A(n2174), .Z(n2181) );
  CIVX2 U3555 ( .A(n2172), .Z(n2182) );
  CIVX2 U3556 ( .A(n2174), .Z(n2184) );
  CIVX2 U3557 ( .A(n2172), .Z(n2186) );
  CIVX2 U3558 ( .A(n2174), .Z(n2187) );
  CIVX2 U3559 ( .A(n2170), .Z(n2189) );
  CIVX2 U3560 ( .A(n2175), .Z(n2190) );
  CIVX2 U3561 ( .A(n2172), .Z(n2191) );
  CIVX2 U3562 ( .A(n2039), .Z(n2192) );
  CIVX2 U3563 ( .A(n2168), .Z(n2193) );
  CIVX2 U3564 ( .A(n2168), .Z(n2194) );
  CIVX2 U3565 ( .A(n2039), .Z(n2195) );
  CIVX2 U3566 ( .A(n2039), .Z(n2196) );
  CIVX2 U3567 ( .A(n2173), .Z(n2199) );
  CIVX2 U3568 ( .A(n2170), .Z(n2201) );
  CMXI2X1 U3569 ( .A0(n5131), .A1(n5132), .S(net78759), .Z(n5158) );
  CND2XL U3570 ( .A(inst_fetch[25]), .B(n1478), .Z(net78759) );
  CND2IXL U3571 ( .B(n3663), .A(n3058), .Z(n3067) );
  CND2IXL U3572 ( .B(n3663), .A(n2846), .Z(n2855) );
  CND2XL U3573 ( .A(N197), .B(n3704), .Z(n2586) );
  CNR2IX1 U3574 ( .B(n2694), .A(n2653), .Z(n2661) );
  CND2X1 U3575 ( .A(n2708), .B(n2709), .Z(N294) );
  CMXI2XL U3576 ( .A0(n2677), .A1(n2676), .S(net87269), .Z(n2678) );
  CNR2XL U3577 ( .A(n2022), .B(net87372), .Z(n2820) );
  CND2XL U3578 ( .A(net87368), .B(n1531), .Z(n3612) );
  CNR2XL U3579 ( .A(n2074), .B(net87389), .Z(n2813) );
  COND1XL U3580 ( .A(net76796), .B(net87691), .C(n5216), .Z(j_type_c) );
  CNR2XL U3581 ( .A(net88116), .B(net87691), .Z(n5215) );
  CMXI2XL U3582 ( .A0(net78792), .A1(net76796), .S(net87691), .Z(n5242) );
  CNR2IXL U3583 ( .B(net87489), .A(n2495), .Z(n2504) );
  CNR2IXL U3584 ( .B(n5227), .A(net88101), .Z(opcode_ext_c[10]) );
  CNR2IXL U3585 ( .B(n5226), .A(net88101), .Z(opcode_ext_c[9]) );
  CNR2IXL U3586 ( .B(n5225), .A(net88101), .Z(opcode_ext_c[8]) );
  CNR2IXL U3587 ( .B(n5224), .A(net88101), .Z(opcode_ext_c[7]) );
  CNR2IXL U3588 ( .B(n5223), .A(net88101), .Z(opcode_ext_c[6]) );
  CNR2IXL U3589 ( .B(n5222), .A(net88101), .Z(opcode_ext_c[5]) );
  CNR2IXL U3590 ( .B(n5221), .A(net88101), .Z(opcode_ext_c[4]) );
  CNR2IXL U3591 ( .B(n5220), .A(net88101), .Z(opcode_ext_c[3]) );
  CNR2IXL U3592 ( .B(n5219), .A(net88101), .Z(opcode_ext_c[2]) );
  CNR2IXL U3593 ( .B(n5218), .A(net88101), .Z(opcode_ext_c[1]) );
  CNR2IXL U3594 ( .B(n5217), .A(net88101), .Z(opcode_ext_c[0]) );
  COND1XL U3595 ( .A(net88101), .B(n5247), .C(n5216), .Z(regc_addr_c[4]) );
  COND1XL U3596 ( .A(net88101), .B(n5248), .C(n5216), .Z(regc_addr_c[3]) );
  COND1XL U3597 ( .A(net88101), .B(n5249), .C(n5216), .Z(regc_addr_c[2]) );
  COND1XL U3598 ( .A(net88101), .B(n5250), .C(n5216), .Z(regc_addr_c[1]) );
  COND1XL U3599 ( .A(net88101), .B(n5251), .C(n5216), .Z(regc_addr_c[0]) );
  CIVX2 U3600 ( .A(net82627), .Z(net82617) );
  CIVX2 U3601 ( .A(net82625), .Z(net82619) );
  CIVX2 U3602 ( .A(net82611), .Z(net82577) );
  CIVX2 U3603 ( .A(net82609), .Z(net82579) );
  CIVX2 U3604 ( .A(net82543), .Z(net82537) );
  CIVX2 U3605 ( .A(net82571), .Z(net82539) );
  CIVX2 U3606 ( .A(net82519), .Z(net82497) );
  CIVX2 U3607 ( .A(net82517), .Z(net82499) );
  CIVX2 U3608 ( .A(net82483), .Z(net82457) );
  CIVX2 U3609 ( .A(net82479), .Z(net82459) );
  CIVX2 U3610 ( .A(net82387), .Z(net82377) );
  CIVX2 U3611 ( .A(net82385), .Z(net82379) );
  CIVX2 U3612 ( .A(n2284), .Z(n2279) );
  CIVX2 U3613 ( .A(n2284), .Z(n2280) );
  CIVX2 U3614 ( .A(n2289), .Z(n2285) );
  CIVX2 U3615 ( .A(n2288), .Z(n2286) );
  CIVX2 U3616 ( .A(n2305), .Z(n2302) );
  CIVX2 U3617 ( .A(n2308), .Z(n2303) );
  CIVX2 U3618 ( .A(n2318), .Z(n2309) );
  CIVX2 U3619 ( .A(n2317), .Z(n2310) );
  CIVX2 U3620 ( .A(n2329), .Z(n2320) );
  CIVX2 U3621 ( .A(n2328), .Z(n2321) );
  CIVX2 U3622 ( .A(n2349), .Z(n2340) );
  CIVX2 U3623 ( .A(n2348), .Z(n2341) );
  CIVX2 U3624 ( .A(n1528), .Z(n2363) );
  CIVX2 U3625 ( .A(n2378), .Z(n2372) );
  CIVX2 U3626 ( .A(n2378), .Z(n2373) );
  CIVX2 U3627 ( .A(n2400), .Z(n2397) );
  CIVX2 U3628 ( .A(n2399), .Z(n2398) );
  CIVX2 U3629 ( .A(n2424), .Z(n2418) );
  CIVX2 U3630 ( .A(n2421), .Z(n2419) );
  CIVX2 U3631 ( .A(n2429), .Z(n2425) );
  CIVX2 U3632 ( .A(n2428), .Z(n2426) );
  CIVX2 U3633 ( .A(n2436), .Z(n2432) );
  CIVX2 U3634 ( .A(n2435), .Z(n2433) );
  CND2X4 U3635 ( .A(r_type), .B(n2455), .Z(n3181) );
  CIVX8 U3636 ( .A(n3181), .Z(n3701) );
  CAOR2X2 U3637 ( .A(data_mem_rdata_i[0]), .B(n2202), .C(alu_op_wb[0]), .D(
        n2207), .Z(n2214) );
  CAOR2X2 U3638 ( .A(data_mem_rdata_i[0]), .B(n2202), .C(alu_op_wb[0]), .D(
        n2206), .Z(n2215) );
  CAOR2X2 U3639 ( .A(data_mem_rdata_i[1]), .B(n2202), .C(alu_op_wb[1]), .D(
        n2207), .Z(n2216) );
  CAOR2X2 U3640 ( .A(data_mem_rdata_i[1]), .B(n2202), .C(alu_op_wb[1]), .D(
        n2205), .Z(n2217) );
  CAOR2X2 U3641 ( .A(data_mem_rdata_i[2]), .B(n2202), .C(alu_op_wb[2]), .D(
        n2209), .Z(net83076) );
  CAOR2X2 U3642 ( .A(data_mem_rdata_i[2]), .B(n2202), .C(alu_op_wb[2]), .D(
        n2208), .Z(net83077) );
  CAOR2X2 U3643 ( .A(data_mem_rdata_i[3]), .B(n2202), .C(alu_op_wb[3]), .D(
        n2213), .Z(n2218) );
  CAOR2X2 U3644 ( .A(data_mem_rdata_i[3]), .B(n2202), .C(alu_op_wb[3]), .D(
        n2212), .Z(n2219) );
  CAOR2X2 U3645 ( .A(data_mem_rdata_i[4]), .B(n2202), .C(alu_op_wb[4]), .D(
        n2205), .Z(net83072) );
  CAOR2X2 U3646 ( .A(data_mem_rdata_i[4]), .B(n2202), .C(alu_op_wb[4]), .D(
        n2204), .Z(net83073) );
  CAOR2X2 U3647 ( .A(data_mem_rdata_i[5]), .B(n2202), .C(alu_op_wb[5]), .D(
        n2209), .Z(n2220) );
  CAOR2X2 U3648 ( .A(data_mem_rdata_i[5]), .B(n2202), .C(alu_op_wb[5]), .D(
        n2208), .Z(n2221) );
  CAOR2X2 U3649 ( .A(data_mem_rdata_i[6]), .B(n2202), .C(alu_op_wb[6]), .D(
        n2210), .Z(n2222) );
  CAOR2X2 U3650 ( .A(data_mem_rdata_i[6]), .B(n2202), .C(alu_op_wb[6]), .D(
        n2206), .Z(n2223) );
  CAOR2X2 U3651 ( .A(data_mem_rdata_i[7]), .B(n2202), .C(alu_op_wb[7]), .D(
        n2212), .Z(n2224) );
  CAOR2X2 U3652 ( .A(data_mem_rdata_i[7]), .B(n2202), .C(alu_op_wb[7]), .D(
        n2211), .Z(n2225) );
  CAOR2X2 U3653 ( .A(data_mem_rdata_i[8]), .B(n2202), .C(alu_op_wb[8]), .D(
        n2207), .Z(n2226) );
  CAOR2X2 U3654 ( .A(data_mem_rdata_i[8]), .B(n2202), .C(alu_op_wb[8]), .D(
        n2206), .Z(n2227) );
  CAOR2X2 U3655 ( .A(data_mem_rdata_i[9]), .B(n2202), .C(alu_op_wb[9]), .D(
        n2209), .Z(n2228) );
  CAOR2X2 U3656 ( .A(data_mem_rdata_i[9]), .B(n2202), .C(alu_op_wb[9]), .D(
        n2208), .Z(n2229) );
  CAOR2X2 U3657 ( .A(data_mem_rdata_i[10]), .B(n2202), .C(alu_op_wb[10]), .D(
        n2211), .Z(n2230) );
  CAOR2X2 U3658 ( .A(data_mem_rdata_i[10]), .B(n2202), .C(alu_op_wb[10]), .D(
        n2210), .Z(n2231) );
  CAOR2X2 U3659 ( .A(data_mem_rdata_i[11]), .B(n2202), .C(alu_op_wb[11]), .D(
        n2213), .Z(net83058) );
  CAOR2X2 U3660 ( .A(data_mem_rdata_i[11]), .B(n2202), .C(alu_op_wb[11]), .D(
        n2207), .Z(net83059) );
  CAOR2X2 U3661 ( .A(data_mem_rdata_i[12]), .B(n2202), .C(alu_op_wb[12]), .D(
        n2205), .Z(n2232) );
  CAOR2X2 U3662 ( .A(data_mem_rdata_i[12]), .B(n2202), .C(alu_op_wb[12]), .D(
        n2204), .Z(n2233) );
  CAOR2X2 U3663 ( .A(data_mem_rdata_i[13]), .B(n2202), .C(alu_op_wb[13]), .D(
        n2211), .Z(net83054) );
  CAOR2X2 U3664 ( .A(data_mem_rdata_i[13]), .B(n2202), .C(alu_op_wb[13]), .D(
        n2210), .Z(net83055) );
  CAOR2X2 U3665 ( .A(data_mem_rdata_i[13]), .B(n2202), .C(alu_op_wb[13]), .D(
        n2212), .Z(n177) );
  CAOR2X2 U3666 ( .A(data_mem_rdata_i[14]), .B(n2202), .C(alu_op_wb[14]), .D(
        n2212), .Z(n2234) );
  CAOR2X2 U3667 ( .A(data_mem_rdata_i[14]), .B(n2202), .C(alu_op_wb[14]), .D(
        n2213), .Z(n2235) );
  CAOR2X2 U3668 ( .A(data_mem_rdata_i[14]), .B(n2202), .C(alu_op_wb[14]), .D(
        n2213), .Z(n176) );
  CAOR2X2 U3669 ( .A(data_mem_rdata_i[15]), .B(n2202), .C(alu_op_wb[15]), .D(
        n2206), .Z(n2236) );
  CAOR2X2 U3670 ( .A(data_mem_rdata_i[15]), .B(n2202), .C(alu_op_wb[15]), .D(
        n2208), .Z(n2237) );
  CAOR2X2 U3671 ( .A(data_mem_rdata_i[15]), .B(n2202), .C(alu_op_wb[15]), .D(
        n2207), .Z(n175) );
  CAOR2X2 U3672 ( .A(data_mem_rdata_i[16]), .B(n2202), .C(alu_op_wb[16]), .D(
        n2204), .Z(n2238) );
  CAOR2X2 U3673 ( .A(data_mem_rdata_i[16]), .B(n2202), .C(alu_op_wb[16]), .D(
        n2208), .Z(n2239) );
  CAOR2X2 U3674 ( .A(data_mem_rdata_i[16]), .B(n2202), .C(alu_op_wb[16]), .D(
        n2205), .Z(n174) );
  CAOR2X2 U3675 ( .A(data_mem_rdata_i[17]), .B(n2202), .C(alu_op_wb[17]), .D(
        n2207), .Z(n2240) );
  CAOR2X2 U3676 ( .A(data_mem_rdata_i[17]), .B(n2202), .C(alu_op_wb[17]), .D(
        n2206), .Z(n2241) );
  CAOR2X2 U3677 ( .A(data_mem_rdata_i[17]), .B(n2202), .C(alu_op_wb[17]), .D(
        n2204), .Z(n173) );
  CAOR2X2 U3678 ( .A(data_mem_rdata_i[18]), .B(n2202), .C(alu_op_wb[18]), .D(
        n2209), .Z(n2242) );
  CAOR2X2 U3679 ( .A(data_mem_rdata_i[18]), .B(n2202), .C(alu_op_wb[18]), .D(
        n2205), .Z(n2243) );
  CAOR2X2 U3680 ( .A(data_mem_rdata_i[18]), .B(n2202), .C(alu_op_wb[18]), .D(
        n2209), .Z(n172) );
  CAOR2X2 U3681 ( .A(data_mem_rdata_i[19]), .B(n2202), .C(alu_op_wb[19]), .D(
        n2211), .Z(n2244) );
  CAOR2X2 U3682 ( .A(data_mem_rdata_i[19]), .B(n2202), .C(alu_op_wb[19]), .D(
        n2210), .Z(n2245) );
  CAOR2X2 U3683 ( .A(data_mem_rdata_i[19]), .B(n2202), .C(alu_op_wb[19]), .D(
        n2208), .Z(n171) );
  CAOR2X2 U3684 ( .A(data_mem_rdata_i[20]), .B(n2202), .C(alu_op_wb[20]), .D(
        n2210), .Z(n2246) );
  CAOR2X2 U3685 ( .A(data_mem_rdata_i[20]), .B(n2202), .C(alu_op_wb[20]), .D(
        n2209), .Z(n2247) );
  CAOR2X2 U3686 ( .A(data_mem_rdata_i[20]), .B(n2202), .C(alu_op_wb[20]), .D(
        n2211), .Z(n170) );
  CAOR2X2 U3687 ( .A(data_mem_rdata_i[21]), .B(n2202), .C(alu_op_wb[21]), .D(
        n2207), .Z(n2248) );
  CAOR2X2 U3688 ( .A(data_mem_rdata_i[21]), .B(n2202), .C(alu_op_wb[21]), .D(
        n2206), .Z(n2249) );
  CAOR2X2 U3689 ( .A(data_mem_rdata_i[21]), .B(n2202), .C(alu_op_wb[21]), .D(
        n2210), .Z(n169) );
  CAOR2X2 U3690 ( .A(data_mem_rdata_i[22]), .B(n2202), .C(alu_op_wb[22]), .D(
        n2213), .Z(n2250) );
  CAOR2X2 U3691 ( .A(data_mem_rdata_i[22]), .B(n2202), .C(alu_op_wb[22]), .D(
        n2212), .Z(n2251) );
  CAOR2X2 U3692 ( .A(data_mem_rdata_i[22]), .B(n2202), .C(alu_op_wb[22]), .D(
        n2204), .Z(n168) );
  CAOR2X2 U3693 ( .A(data_mem_rdata_i[23]), .B(n2202), .C(alu_op_wb[23]), .D(
        n2213), .Z(n2252) );
  CAOR2X2 U3694 ( .A(data_mem_rdata_i[23]), .B(n2202), .C(alu_op_wb[23]), .D(
        n2212), .Z(n2253) );
  CAOR2X2 U3695 ( .A(data_mem_rdata_i[23]), .B(n2202), .C(alu_op_wb[23]), .D(
        n2204), .Z(n167) );
  CAOR2X2 U3696 ( .A(data_mem_rdata_i[24]), .B(n2202), .C(alu_op_wb[24]), .D(
        n2208), .Z(n2254) );
  CAOR2X2 U3697 ( .A(data_mem_rdata_i[24]), .B(n2202), .C(alu_op_wb[24]), .D(
        n2205), .Z(n2255) );
  CAOR2X2 U3698 ( .A(data_mem_rdata_i[24]), .B(n2202), .C(alu_op_wb[24]), .D(
        n2209), .Z(n166) );
  CAOR2X2 U3699 ( .A(data_mem_rdata_i[25]), .B(n2202), .C(alu_op_wb[25]), .D(
        n2205), .Z(n2256) );
  CAOR2X2 U3700 ( .A(data_mem_rdata_i[25]), .B(n2202), .C(alu_op_wb[25]), .D(
        n2211), .Z(n2257) );
  CAOR2X2 U3701 ( .A(data_mem_rdata_i[25]), .B(n2202), .C(alu_op_wb[25]), .D(
        n2206), .Z(n165) );
  CAOR2X2 U3702 ( .A(data_mem_rdata_i[26]), .B(n2202), .C(alu_op_wb[26]), .D(
        n2206), .Z(n2258) );
  CAOR2X2 U3703 ( .A(data_mem_rdata_i[26]), .B(n2202), .C(alu_op_wb[26]), .D(
        n2207), .Z(n2259) );
  CAOR2X2 U3704 ( .A(data_mem_rdata_i[26]), .B(n2202), .C(alu_op_wb[26]), .D(
        n2207), .Z(n164) );
  CAOR2X2 U3705 ( .A(data_mem_rdata_i[27]), .B(n2202), .C(alu_op_wb[27]), .D(
        n2209), .Z(n2260) );
  CAOR2X2 U3706 ( .A(data_mem_rdata_i[27]), .B(n2202), .C(alu_op_wb[27]), .D(
        n2208), .Z(n2261) );
  CAOR2X2 U3707 ( .A(data_mem_rdata_i[27]), .B(n2202), .C(alu_op_wb[27]), .D(
        n2210), .Z(n163) );
  CAOR2X2 U3708 ( .A(data_mem_rdata_i[28]), .B(n2202), .C(alu_op_wb[28]), .D(
        n2212), .Z(n2262) );
  CAOR2X2 U3709 ( .A(data_mem_rdata_i[28]), .B(n2202), .C(alu_op_wb[28]), .D(
        n2211), .Z(n2263) );
  CAOR2X2 U3710 ( .A(data_mem_rdata_i[28]), .B(n2202), .C(alu_op_wb[28]), .D(
        n2208), .Z(n162) );
  CAOR2X2 U3711 ( .A(data_mem_rdata_i[29]), .B(n2202), .C(alu_op_wb[29]), .D(
        n2210), .Z(n2264) );
  CAOR2X2 U3712 ( .A(data_mem_rdata_i[29]), .B(n2202), .C(alu_op_wb[29]), .D(
        n2209), .Z(n2265) );
  CAOR2X2 U3713 ( .A(data_mem_rdata_i[29]), .B(n2202), .C(alu_op_wb[29]), .D(
        n2210), .Z(n161) );
  CAOR2X2 U3714 ( .A(data_mem_rdata_i[30]), .B(n2202), .C(alu_op_wb[30]), .D(
        n2212), .Z(n2266) );
  CAOR2X2 U3715 ( .A(data_mem_rdata_i[30]), .B(n2202), .C(alu_op_wb[30]), .D(
        n2211), .Z(n2267) );
  CAOR2X2 U3716 ( .A(data_mem_rdata_i[30]), .B(n2202), .C(alu_op_wb[30]), .D(
        n2213), .Z(n160) );
  CAOR2X2 U3717 ( .A(data_mem_rdata_i[31]), .B(data_mem_rd_d), .C(
        alu_op_wb[31]), .D(n2213), .Z(n2268) );
  CAOR2X2 U3718 ( .A(data_mem_rdata_i[31]), .B(data_mem_rd_d), .C(
        alu_op_wb[31]), .D(n2212), .Z(n2269) );
  CIVXL U3719 ( .A(n238), .Z(net82665) );
  CIVXL U3720 ( .A(n238), .Z(net82667) );
  CIVXL U3721 ( .A(n238), .Z(net82677) );
  CIVXL U3722 ( .A(n238), .Z(net82679) );
  CIVXL U3723 ( .A(n238), .Z(net82683) );
  CIVXL U3724 ( .A(n238), .Z(net82689) );
  CIVXL U3725 ( .A(net82643), .Z(net82621) );
  CIVXL U3726 ( .A(n237), .Z(net82625) );
  CIVXL U3727 ( .A(n237), .Z(net82627) );
  CIVXL U3728 ( .A(n237), .Z(net82639) );
  CIVXL U3729 ( .A(n237), .Z(net82643) );
  CIVXL U3730 ( .A(net82583), .Z(net82581) );
  CIVXL U3731 ( .A(n236), .Z(net82583) );
  CIVXL U3732 ( .A(n236), .Z(net82585) );
  CIVXL U3733 ( .A(n236), .Z(net82587) );
  CIVXL U3734 ( .A(n236), .Z(net82591) );
  CIVXL U3735 ( .A(n236), .Z(net82593) );
  CIVXL U3736 ( .A(n236), .Z(net82597) );
  CIVXL U3737 ( .A(n236), .Z(net82599) );
  CIVXL U3738 ( .A(n236), .Z(net82603) );
  CIVXL U3739 ( .A(n236), .Z(net82605) );
  CIVXL U3740 ( .A(n236), .Z(net82609) );
  CIVXL U3741 ( .A(n236), .Z(net82611) );
  CIVXL U3742 ( .A(net82557), .Z(net82541) );
  CIVXL U3743 ( .A(n235), .Z(net82543) );
  CIVXL U3744 ( .A(n235), .Z(net82549) );
  CIVXL U3745 ( .A(n235), .Z(net82557) );
  CIVXL U3746 ( .A(n235), .Z(net82571) );
  CIVXL U3747 ( .A(net82503), .Z(net82501) );
  CIVXL U3748 ( .A(n234), .Z(net82503) );
  CIVXL U3749 ( .A(n234), .Z(net82505) );
  CIVXL U3750 ( .A(n234), .Z(net82507) );
  CIVXL U3751 ( .A(n234), .Z(net82509) );
  CIVXL U3752 ( .A(n234), .Z(net82513) );
  CIVXL U3753 ( .A(n234), .Z(net82515) );
  CIVXL U3754 ( .A(n234), .Z(net82517) );
  CIVXL U3755 ( .A(n234), .Z(net82519) );
  CIVXL U3756 ( .A(n234), .Z(net82521) );
  CIVXL U3757 ( .A(n234), .Z(net82523) );
  CIVXL U3758 ( .A(n234), .Z(net82527) );
  CIVXL U3759 ( .A(n234), .Z(net82529) );
  CIVXL U3760 ( .A(n234), .Z(net82533) );
  CIVXL U3761 ( .A(net82485), .Z(net82461) );
  CIVXL U3762 ( .A(n233), .Z(net82463) );
  CIVXL U3763 ( .A(n233), .Z(net82465) );
  CIVXL U3764 ( .A(n233), .Z(net82469) );
  CIVXL U3765 ( .A(n233), .Z(net82473) );
  CIVXL U3766 ( .A(n233), .Z(net82477) );
  CIVXL U3767 ( .A(n233), .Z(net82479) );
  CIVXL U3768 ( .A(n233), .Z(net82483) );
  CIVXL U3769 ( .A(n233), .Z(net82485) );
  CIVXL U3770 ( .A(n233), .Z(net82489) );
  CIVXL U3771 ( .A(n233), .Z(net82491) );
  CIVXL U3772 ( .A(net87043), .Z(net82421) );
  CIVXL U3773 ( .A(net87042), .Z(net82425) );
  CIVXL U3774 ( .A(net87042), .Z(net82427) );
  CIVXL U3775 ( .A(net87042), .Z(net82437) );
  CIVXL U3776 ( .A(net87042), .Z(net82439) );
  CIVXL U3777 ( .A(net87042), .Z(net82443) );
  CIVXL U3778 ( .A(net82403), .Z(net82381) );
  CIVXL U3779 ( .A(n227), .Z(net82385) );
  CIVXL U3780 ( .A(n227), .Z(net82387) );
  CIVXL U3781 ( .A(n227), .Z(net82399) );
  CIVXL U3782 ( .A(n227), .Z(net82403) );
  CIVXL U3783 ( .A(n226), .Z(n2281) );
  CIVXL U3784 ( .A(n226), .Z(n2282) );
  CIVXL U3785 ( .A(n226), .Z(n2283) );
  CIVXL U3786 ( .A(n226), .Z(n2284) );
  CIVXL U3787 ( .A(n2291), .Z(n2287) );
  CIVXL U3788 ( .A(n225), .Z(n2288) );
  CIVXL U3789 ( .A(n225), .Z(n2289) );
  CIVXL U3790 ( .A(n225), .Z(n2290) );
  CIVXL U3791 ( .A(n225), .Z(n2291) );
  CIVXL U3792 ( .A(n224), .Z(n2292) );
  CIVXL U3793 ( .A(n224), .Z(n2293) );
  CIVXL U3794 ( .A(n224), .Z(n2294) );
  CIVXL U3795 ( .A(n224), .Z(n2295) );
  CIVXL U3796 ( .A(n224), .Z(n2296) );
  CIVXL U3797 ( .A(n224), .Z(n2297) );
  CIVXL U3798 ( .A(n224), .Z(n2298) );
  CIVXL U3799 ( .A(n224), .Z(n2299) );
  CIVXL U3800 ( .A(n224), .Z(n2300) );
  CIVXL U3801 ( .A(n224), .Z(n2301) );
  CIVXL U3802 ( .A(n2307), .Z(n2304) );
  CIVXL U3803 ( .A(n223), .Z(n2305) );
  CIVXL U3804 ( .A(n223), .Z(n2306) );
  CIVXL U3805 ( .A(n223), .Z(n2307) );
  CIVXL U3806 ( .A(n223), .Z(n2308) );
  CIVXL U3807 ( .A(n2319), .Z(n2311) );
  CIVXL U3808 ( .A(n222), .Z(n2312) );
  CIVXL U3809 ( .A(n222), .Z(n2313) );
  CIVXL U3810 ( .A(n222), .Z(n2314) );
  CIVXL U3811 ( .A(n222), .Z(n2315) );
  CIVXL U3812 ( .A(n222), .Z(n2316) );
  CIVXL U3813 ( .A(n222), .Z(n2317) );
  CIVXL U3814 ( .A(n222), .Z(n2318) );
  CIVXL U3815 ( .A(n222), .Z(n2319) );
  CIVXL U3816 ( .A(n2330), .Z(n2322) );
  CIVXL U3817 ( .A(n221), .Z(n2323) );
  CIVXL U3818 ( .A(n221), .Z(n2324) );
  CIVXL U3819 ( .A(n221), .Z(n2325) );
  CIVXL U3820 ( .A(n221), .Z(n2326) );
  CIVXL U3821 ( .A(n221), .Z(n2327) );
  CIVXL U3822 ( .A(n221), .Z(n2328) );
  CIVXL U3823 ( .A(n221), .Z(n2329) );
  CIVXL U3824 ( .A(n221), .Z(n2330) );
  CIVXL U3825 ( .A(n1526), .Z(n2331) );
  CIVXL U3826 ( .A(n220), .Z(n2332) );
  CIVXL U3827 ( .A(n220), .Z(n2333) );
  CIVXL U3828 ( .A(n220), .Z(n2334) );
  CIVXL U3829 ( .A(n220), .Z(n2335) );
  CIVXL U3830 ( .A(n220), .Z(n2336) );
  CIVXL U3831 ( .A(n220), .Z(n2337) );
  CIVXL U3832 ( .A(n220), .Z(n2338) );
  CIVXL U3833 ( .A(n220), .Z(n2339) );
  CIVXL U3834 ( .A(n2350), .Z(n2342) );
  CIVXL U3835 ( .A(n218), .Z(n2343) );
  CIVXL U3836 ( .A(n218), .Z(n2344) );
  CIVXL U3837 ( .A(n218), .Z(n2345) );
  CIVXL U3838 ( .A(n218), .Z(n2346) );
  CIVXL U3839 ( .A(n218), .Z(n2347) );
  CIVXL U3840 ( .A(n218), .Z(n2348) );
  CIVXL U3841 ( .A(n218), .Z(n2349) );
  CIVXL U3842 ( .A(n218), .Z(n2350) );
  CIVXL U3843 ( .A(net82051), .Z(net82021) );
  CIVXL U3844 ( .A(n217), .Z(net82025) );
  CIVXL U3845 ( .A(n217), .Z(net82027) );
  CIVXL U3846 ( .A(n217), .Z(net82031) );
  CIVXL U3847 ( .A(n217), .Z(net82037) );
  CIVXL U3848 ( .A(n217), .Z(net82039) );
  CIVXL U3849 ( .A(n217), .Z(net82043) );
  CIVXL U3850 ( .A(n217), .Z(net82051) );
  CIVXL U3851 ( .A(net82011), .Z(net81981) );
  CIVXL U3852 ( .A(n216), .Z(net81985) );
  CIVXL U3853 ( .A(n216), .Z(net81987) );
  CIVXL U3854 ( .A(n216), .Z(net81991) );
  CIVXL U3855 ( .A(n216), .Z(net81997) );
  CIVXL U3856 ( .A(n216), .Z(net81999) );
  CIVXL U3857 ( .A(n216), .Z(net82011) );
  CIVXL U3858 ( .A(net81971), .Z(net81941) );
  CIVXL U3859 ( .A(n215), .Z(net81945) );
  CIVXL U3860 ( .A(n215), .Z(net81947) );
  CIVXL U3861 ( .A(n215), .Z(net81951) );
  CIVXL U3862 ( .A(n215), .Z(net81957) );
  CIVXL U3863 ( .A(n215), .Z(net81959) );
  CIVXL U3864 ( .A(n215), .Z(net81971) );
  CIVXL U3865 ( .A(n1516), .Z(net81901) );
  CIVXL U3866 ( .A(n214), .Z(net81905) );
  CIVXL U3867 ( .A(n214), .Z(net81907) );
  CIVXL U3868 ( .A(n214), .Z(net81917) );
  CIVXL U3869 ( .A(n214), .Z(net81919) );
  CIVXL U3870 ( .A(n214), .Z(net81923) );
  CIVXL U3871 ( .A(n1518), .Z(n2351) );
  CIVXL U3872 ( .A(n213), .Z(n2352) );
  CIVXL U3873 ( .A(n213), .Z(n2353) );
  CIVXL U3874 ( .A(n213), .Z(n2354) );
  CIVXL U3875 ( .A(n213), .Z(n2355) );
  CIVXL U3876 ( .A(n213), .Z(n2356) );
  CIVXL U3877 ( .A(n1520), .Z(n2357) );
  CIVXL U3878 ( .A(n212), .Z(n2358) );
  CIVXL U3879 ( .A(n212), .Z(n2359) );
  CIVXL U3880 ( .A(n212), .Z(n2360) );
  CIVXL U3881 ( .A(n212), .Z(n2361) );
  CIVXL U3882 ( .A(n212), .Z(n2362) );
  CIVXL U3883 ( .A(n211), .Z(n2364) );
  CIVXL U3884 ( .A(n211), .Z(n2365) );
  CIVXL U3885 ( .A(n211), .Z(n2366) );
  CIVXL U3886 ( .A(n211), .Z(n2367) );
  CIVXL U3887 ( .A(n211), .Z(n2368) );
  CIVXL U3888 ( .A(n211), .Z(n2369) );
  CIVXL U3889 ( .A(n211), .Z(n2370) );
  CIVXL U3890 ( .A(n211), .Z(n2371) );
  CIVXL U3891 ( .A(n2378), .Z(n2374) );
  CIVXL U3892 ( .A(n1940), .Z(n2375) );
  CIVXL U3893 ( .A(n1940), .Z(n2376) );
  CIVXL U3894 ( .A(n1940), .Z(n2377) );
  CIVXL U3895 ( .A(n209), .Z(n2378) );
  CIVXL U3896 ( .A(n2382), .Z(n2379) );
  CIVXL U3897 ( .A(n205), .Z(n2380) );
  CIVXL U3898 ( .A(n205), .Z(n2381) );
  CIVXL U3899 ( .A(n205), .Z(n2382) );
  CIVXL U3900 ( .A(n205), .Z(n2383) );
  CIVXL U3901 ( .A(n205), .Z(n2384) );
  CIVXL U3902 ( .A(n205), .Z(n2385) );
  CIVXL U3903 ( .A(n205), .Z(n2386) );
  CIVXL U3904 ( .A(n205), .Z(n2387) );
  CIVXL U3905 ( .A(n2391), .Z(n2388) );
  CIVXL U3906 ( .A(n203), .Z(n2389) );
  CIVXL U3907 ( .A(n203), .Z(n2390) );
  CIVXL U3908 ( .A(n203), .Z(n2391) );
  CIVXL U3909 ( .A(n203), .Z(n2392) );
  CIVXL U3910 ( .A(n203), .Z(n2393) );
  CIVXL U3911 ( .A(n203), .Z(n2394) );
  CIVXL U3912 ( .A(n203), .Z(n2395) );
  CIVXL U3913 ( .A(n203), .Z(n2396) );
  CIVXL U3914 ( .A(n201), .Z(n2399) );
  CIVXL U3915 ( .A(n201), .Z(n2400) );
  CIVXL U3916 ( .A(n201), .Z(n2401) );
  CIVXL U3917 ( .A(n201), .Z(n2402) );
  CIVXL U3918 ( .A(n2404), .Z(n2403) );
  CIVXL U3919 ( .A(n199), .Z(n2405) );
  CIVXL U3920 ( .A(n199), .Z(n2406) );
  CIVXL U3921 ( .A(n199), .Z(n2407) );
  CIVXL U3922 ( .A(n199), .Z(n2408) );
  CIVXL U3923 ( .A(n2410), .Z(n2409) );
  CIVXL U3924 ( .A(n197), .Z(n2411) );
  CIVXL U3925 ( .A(n197), .Z(n2412) );
  CIVXL U3926 ( .A(n197), .Z(n2413) );
  CIVXL U3927 ( .A(n197), .Z(n2414) );
  CIVXL U3928 ( .A(n197), .Z(n2415) );
  CIVXL U3929 ( .A(n197), .Z(n2416) );
  CIVXL U3930 ( .A(n197), .Z(n2417) );
  CIVXL U3931 ( .A(n2423), .Z(n2420) );
  CIVXL U3932 ( .A(n195), .Z(n2421) );
  CIVXL U3933 ( .A(n195), .Z(n2422) );
  CIVXL U3934 ( .A(n195), .Z(n2423) );
  CIVXL U3935 ( .A(n195), .Z(n2424) );
  CIVXL U3936 ( .A(n2431), .Z(n2427) );
  CIVXL U3937 ( .A(n193), .Z(n2428) );
  CIVXL U3938 ( .A(n193), .Z(n2429) );
  CIVXL U3939 ( .A(n193), .Z(n2430) );
  CIVXL U3940 ( .A(n2438), .Z(n2434) );
  CIVXL U3941 ( .A(n158), .Z(n2435) );
  CIVXL U3942 ( .A(n158), .Z(n2436) );
  CIVXL U3943 ( .A(n158), .Z(n2437) );
  CIVXL U3944 ( .A(n158), .Z(n2438) );
  CIVX2 U3945 ( .A(immi_val[31]), .Z(n5246) );
  CND2IX1 U3946 ( .B(opcode_ex[5]), .A(opcode_ex[2]), .Z(n2439) );
  CIVX2 U3947 ( .A(n2439), .Z(n5239) );
  CND2X2 U3948 ( .A(n2440), .B(n2156), .Z(n2443) );
  CIVX2 U3949 ( .A(n2443), .Z(n2441) );
  CIVX2 U3950 ( .A(n338), .Z(n2447) );
  CND2IX1 U3951 ( .B(opcode_ex[0]), .A(opcode_ex[1]), .Z(n2442) );
  CIVX2 U3952 ( .A(n2442), .Z(n2449) );
  CND3X2 U3953 ( .A(opcode_ex[3]), .B(opcode_ex[4]), .C(n2449), .Z(n3332) );
  CIVX2 U3954 ( .A(opcode_ex[2]), .Z(n2445) );
  CIVX2 U3955 ( .A(opcode_ex[5]), .Z(n5240) );
  CNR2IX2 U3956 ( .B(n5240), .A(n2443), .Z(n2444) );
  CND2X2 U3957 ( .A(n2445), .B(n2444), .Z(n3699) );
  CIVX2 U3958 ( .A(n3699), .Z(n3476) );
  CND2X2 U3959 ( .A(n2447), .B(n2446), .Z(n2455) );
  CIVX2 U3960 ( .A(opcode_ex[4]), .Z(n2454) );
  COND3X1 U3961 ( .A(n5239), .B(n2454), .C(n2450), .D(n2449), .Z(n2451) );
  CND2X2 U3962 ( .A(N31), .B(n2147), .Z(n3330) );
  CND2X2 U3963 ( .A(n2135), .B(n3330), .Z(n3344) );
  CMXI2X1 U3964 ( .A0(\reg_mem[0][0] ), .A1(\reg_mem[1][0] ), .S(net87396), 
        .Z(n2463) );
  CMXI2X1 U3965 ( .A0(\reg_mem[2][0] ), .A1(\reg_mem[3][0] ), .S(net87389), 
        .Z(n2462) );
  CMXI2X1 U3966 ( .A0(n2463), .A1(n2462), .S(n2179), .Z(n2467) );
  CMXI2X1 U3967 ( .A0(\reg_mem[4][0] ), .A1(\reg_mem[5][0] ), .S(net87392), 
        .Z(n2465) );
  CMXI2X1 U3968 ( .A0(\reg_mem[6][0] ), .A1(\reg_mem[7][0] ), .S(net87411), 
        .Z(n2464) );
  CMXI2X1 U3969 ( .A0(n2465), .A1(n2464), .S(n2185), .Z(n2466) );
  CMXI2X1 U3970 ( .A0(n2467), .A1(n2466), .S(net87279), .Z(n2475) );
  CMXI2X1 U3971 ( .A0(\reg_mem[8][0] ), .A1(\reg_mem[9][0] ), .S(net87386), 
        .Z(n2469) );
  CMXI2X1 U3972 ( .A0(\reg_mem[10][0] ), .A1(\reg_mem[11][0] ), .S(net87392), 
        .Z(n2468) );
  CMXI2X1 U3973 ( .A0(n2469), .A1(n2468), .S(n2180), .Z(n2473) );
  CMXI2X1 U3974 ( .A0(\reg_mem[14][0] ), .A1(\reg_mem[15][0] ), .S(net87386), 
        .Z(n2470) );
  CMXI2X1 U3975 ( .A0(n2471), .A1(n2470), .S(n2165), .Z(n2472) );
  CMXI2X1 U3976 ( .A0(n2473), .A1(n2472), .S(net87255), .Z(n2474) );
  CMXI2X1 U3977 ( .A0(n2475), .A1(n2474), .S(n1532), .Z(n2491) );
  CMXI2X1 U3978 ( .A0(\reg_mem[16][0] ), .A1(\reg_mem[17][0] ), .S(net87409), 
        .Z(n2477) );
  CMXI2X1 U3979 ( .A0(\reg_mem[18][0] ), .A1(\reg_mem[19][0] ), .S(net87411), 
        .Z(n2476) );
  CMXI2X1 U3980 ( .A0(n2477), .A1(n2476), .S(n2186), .Z(n2481) );
  CMXI2X1 U3981 ( .A0(\reg_mem[20][0] ), .A1(\reg_mem[21][0] ), .S(net87395), 
        .Z(n2479) );
  CMXI2X1 U3982 ( .A0(\reg_mem[22][0] ), .A1(\reg_mem[23][0] ), .S(net87385), 
        .Z(n2478) );
  CMXI2X1 U3983 ( .A0(n2479), .A1(n2478), .S(n2190), .Z(n2480) );
  CMXI2X1 U3984 ( .A0(\reg_mem[24][0] ), .A1(\reg_mem[25][0] ), .S(net87396), 
        .Z(n2483) );
  CMXI2X1 U3985 ( .A0(\reg_mem[26][0] ), .A1(\reg_mem[27][0] ), .S(net87397), 
        .Z(n2482) );
  CMXI2X1 U3986 ( .A0(n2483), .A1(n2482), .S(n2166), .Z(n2487) );
  CMXI2X1 U3987 ( .A0(\reg_mem[28][0] ), .A1(\reg_mem[29][0] ), .S(net87405), 
        .Z(n2485) );
  CMXI2X1 U3988 ( .A0(\reg_mem[30][0] ), .A1(\reg_mem[31][0] ), .S(net87395), 
        .Z(n2484) );
  CMXI2X1 U3989 ( .A0(n2485), .A1(n2484), .S(n2191), .Z(n2486) );
  CMXI2X1 U3990 ( .A0(n2487), .A1(n2486), .S(net87258), .Z(n2488) );
  CIVX2 U3991 ( .A(alu_op_c[0]), .Z(n2505) );
  CMXI2X1 U3992 ( .A0(n2494), .A1(inst_fetch[27]), .S(regb_addr[0]), .Z(n2495)
         );
  CMXI2X1 U3993 ( .A0(\reg_mem[0][29] ), .A1(\reg_mem[16][29] ), .S(n2101), 
        .Z(n2508) );
  CMXI2X1 U3994 ( .A0(\reg_mem[6][29] ), .A1(\reg_mem[22][29] ), .S(n2095), 
        .Z(n2509) );
  CMXI2X1 U3995 ( .A0(\reg_mem[8][29] ), .A1(\reg_mem[24][29] ), .S(n2088), 
        .Z(n2514) );
  CMXI2X1 U3996 ( .A0(\reg_mem[10][29] ), .A1(\reg_mem[26][29] ), .S(n2082), 
        .Z(n2513) );
  CMXI2X1 U3997 ( .A0(\reg_mem[12][29] ), .A1(\reg_mem[28][29] ), .S(n2093), 
        .Z(n2516) );
  CMXI2X1 U3998 ( .A0(\reg_mem[14][29] ), .A1(\reg_mem[30][29] ), .S(n2085), 
        .Z(n2515) );
  CMXI2X1 U3999 ( .A0(n2516), .A1(n2515), .S(n2179), .Z(n2517) );
  CMXI2X1 U4000 ( .A0(\reg_mem[1][29] ), .A1(\reg_mem[17][29] ), .S(n2098), 
        .Z(n2522) );
  CMXI2X1 U4001 ( .A0(\reg_mem[5][29] ), .A1(\reg_mem[21][29] ), .S(n1975), 
        .Z(n2524) );
  CMXI2X1 U4002 ( .A0(\reg_mem[7][29] ), .A1(\reg_mem[23][29] ), .S(n2091), 
        .Z(n2523) );
  CMXI2X1 U4003 ( .A0(n2524), .A1(n2523), .S(n2194), .Z(n2525) );
  CMXI2X1 U4004 ( .A0(\reg_mem[9][29] ), .A1(\reg_mem[25][29] ), .S(n1975), 
        .Z(n2528) );
  CMXI2X1 U4005 ( .A0(n2528), .A1(n2527), .S(n2177), .Z(n2532) );
  CMXI2X1 U4006 ( .A0(\reg_mem[13][29] ), .A1(\reg_mem[29][29] ), .S(n2100), 
        .Z(n2530) );
  CMXI2X1 U4007 ( .A0(\reg_mem[15][29] ), .A1(\reg_mem[31][29] ), .S(n2082), 
        .Z(n2529) );
  CMXI2X1 U4008 ( .A0(n2530), .A1(n2529), .S(n2181), .Z(n2531) );
  CMXI2X1 U4009 ( .A0(n2532), .A1(n2531), .S(net87279), .Z(n2533) );
  CIVX2 U4010 ( .A(N125), .Z(n2538) );
  CND2IX1 U4011 ( .B(n3181), .A(N166), .Z(n2540) );
  CND2IX1 U4012 ( .B(n2545), .A(n2544), .Z(alu_op_c[29]) );
  CMXI2X1 U4013 ( .A0(\reg_mem[9][28] ), .A1(\reg_mem[25][28] ), .S(n2093), 
        .Z(n2547) );
  CMXI2X1 U4014 ( .A0(\reg_mem[11][28] ), .A1(\reg_mem[27][28] ), .S(n2088), 
        .Z(n2546) );
  CMXI2X1 U4015 ( .A0(n2547), .A1(n2546), .S(n2165), .Z(n2551) );
  CMXI2X1 U4016 ( .A0(\reg_mem[13][28] ), .A1(\reg_mem[29][28] ), .S(n2095), 
        .Z(n2549) );
  CMXI2X1 U4017 ( .A0(\reg_mem[15][28] ), .A1(\reg_mem[31][28] ), .S(n2100), 
        .Z(n2548) );
  CMXI2X1 U4018 ( .A0(n2549), .A1(n2548), .S(n2189), .Z(n2550) );
  CMXI2X1 U4019 ( .A0(n2551), .A1(n2550), .S(net87278), .Z(n2552) );
  CND2IX1 U4020 ( .B(n3604), .A(n2552), .Z(n2561) );
  CMXI2X1 U4021 ( .A0(\reg_mem[2][28] ), .A1(\reg_mem[18][28] ), .S(n2092), 
        .Z(n2553) );
  CMXI2X1 U4022 ( .A0(n2554), .A1(n2553), .S(n1469), .Z(n2558) );
  CMXI2X1 U4023 ( .A0(\reg_mem[6][28] ), .A1(\reg_mem[22][28] ), .S(n2100), 
        .Z(n2555) );
  CMXI2X1 U4024 ( .A0(n2558), .A1(n2557), .S(n1480), .Z(n2559) );
  CND2IX1 U4025 ( .B(n3612), .A(n2559), .Z(n2560) );
  CMXI2X1 U4026 ( .A0(\reg_mem[8][28] ), .A1(\reg_mem[24][28] ), .S(n2084), 
        .Z(n2563) );
  CMXI2X1 U4027 ( .A0(\reg_mem[10][28] ), .A1(\reg_mem[26][28] ), .S(n2094), 
        .Z(n2562) );
  CMXI2X1 U4028 ( .A0(n2563), .A1(n2562), .S(n2195), .Z(n2567) );
  CMXI2X1 U4029 ( .A0(\reg_mem[12][28] ), .A1(\reg_mem[28][28] ), .S(n2087), 
        .Z(n2565) );
  CMXI2X1 U4030 ( .A0(\reg_mem[14][28] ), .A1(\reg_mem[30][28] ), .S(n2082), 
        .Z(n2564) );
  CMXI2X1 U4031 ( .A0(n2565), .A1(n2564), .S(n2197), .Z(n2566) );
  CMXI2X1 U4032 ( .A0(n2567), .A1(n2566), .S(net87268), .Z(n2568) );
  CMXI2X1 U4033 ( .A0(\reg_mem[1][28] ), .A1(\reg_mem[17][28] ), .S(n2093), 
        .Z(n2570) );
  CMXI2X1 U4034 ( .A0(\reg_mem[3][28] ), .A1(\reg_mem[19][28] ), .S(n1975), 
        .Z(n2569) );
  CMXI2X1 U4035 ( .A0(\reg_mem[5][28] ), .A1(\reg_mem[21][28] ), .S(n2100), 
        .Z(n2572) );
  CMXI2X1 U4036 ( .A0(\reg_mem[7][28] ), .A1(\reg_mem[23][28] ), .S(n2095), 
        .Z(n2571) );
  CMXI2X1 U4037 ( .A0(n2572), .A1(n2571), .S(n2186), .Z(n2573) );
  CMXI2X1 U4038 ( .A0(n2574), .A1(n2573), .S(net87272), .Z(n2575) );
  CND2IX1 U4039 ( .B(n3631), .A(n2575), .Z(n2576) );
  CIVX2 U4040 ( .A(N124), .Z(n2578) );
  CMXI2X1 U4041 ( .A0(\reg_mem[9][27] ), .A1(\reg_mem[25][27] ), .S(n2101), 
        .Z(n2589) );
  CMXI2X1 U4042 ( .A0(\reg_mem[11][27] ), .A1(\reg_mem[27][27] ), .S(n2097), 
        .Z(n2588) );
  CMXI2X1 U4043 ( .A0(n2589), .A1(n2588), .S(n2176), .Z(n2593) );
  CMXI2X1 U4044 ( .A0(\reg_mem[15][27] ), .A1(\reg_mem[31][27] ), .S(n2099), 
        .Z(n2590) );
  CMXI2X1 U4045 ( .A0(n2591), .A1(n2590), .S(n2166), .Z(n2592) );
  CMXI2X1 U4046 ( .A0(n2593), .A1(n2592), .S(net87265), .Z(n2594) );
  CND2IX1 U4047 ( .B(n3604), .A(n2594), .Z(n2603) );
  CMXI2X1 U4048 ( .A0(\reg_mem[2][27] ), .A1(\reg_mem[18][27] ), .S(n2092), 
        .Z(n2595) );
  CMXI2X1 U4049 ( .A0(n2596), .A1(n2595), .S(n2180), .Z(n2600) );
  CMXI2X1 U4050 ( .A0(\reg_mem[4][27] ), .A1(\reg_mem[20][27] ), .S(n2098), 
        .Z(n2598) );
  CMXI2X1 U4051 ( .A0(\reg_mem[6][27] ), .A1(\reg_mem[22][27] ), .S(n2094), 
        .Z(n2597) );
  CMXI2X1 U4052 ( .A0(n2598), .A1(n2597), .S(n2192), .Z(n2599) );
  CMXI2X1 U4053 ( .A0(n2600), .A1(n2599), .S(net87262), .Z(n2601) );
  CND2IX1 U4054 ( .B(n3612), .A(n2601), .Z(n2602) );
  CMXI2X1 U4055 ( .A0(\reg_mem[8][27] ), .A1(\reg_mem[24][27] ), .S(n2097), 
        .Z(n2605) );
  CMXI2X1 U4056 ( .A0(\reg_mem[12][27] ), .A1(\reg_mem[28][27] ), .S(n2104), 
        .Z(n2607) );
  CMXI2X1 U4057 ( .A0(\reg_mem[14][27] ), .A1(\reg_mem[30][27] ), .S(n2097), 
        .Z(n2606) );
  CMXI2X1 U4058 ( .A0(n2607), .A1(n2606), .S(n2196), .Z(n2608) );
  CMXI2X1 U4059 ( .A0(n2609), .A1(n2608), .S(net87273), .Z(n2610) );
  CND2IX1 U4060 ( .B(n3623), .A(n2610), .Z(n2619) );
  CMXI2X1 U4061 ( .A0(\reg_mem[1][27] ), .A1(\reg_mem[17][27] ), .S(n2102), 
        .Z(n2612) );
  CMXI2X1 U4062 ( .A0(\reg_mem[3][27] ), .A1(\reg_mem[19][27] ), .S(n2104), 
        .Z(n2611) );
  CMXI2X1 U4063 ( .A0(n2612), .A1(n2611), .S(n2183), .Z(n2616) );
  CMXI2X1 U4064 ( .A0(\reg_mem[7][27] ), .A1(\reg_mem[23][27] ), .S(n2098), 
        .Z(n2613) );
  CMXI2X1 U4065 ( .A0(n2614), .A1(n2613), .S(n2185), .Z(n2615) );
  CMXI2X1 U4066 ( .A0(n2616), .A1(n2615), .S(net87269), .Z(n2617) );
  CND2IX1 U4067 ( .B(n3631), .A(n2617), .Z(n2618) );
  CIVX2 U4068 ( .A(N123), .Z(n2620) );
  CND2IX1 U4069 ( .B(n2629), .A(n2628), .Z(alu_op_c[27]) );
  CIVX2 U4070 ( .A(\reg_mem[9][26] ), .Z(n4935) );
  CIVX2 U4071 ( .A(\reg_mem[25][26] ), .Z(n4965) );
  CMXI2X1 U4072 ( .A0(n4935), .A1(n4965), .S(n2102), .Z(n2634) );
  CIVX2 U4073 ( .A(\reg_mem[11][26] ), .Z(n4937) );
  CIVX2 U4074 ( .A(\reg_mem[27][26] ), .Z(n4967) );
  CIVX2 U4075 ( .A(\reg_mem[13][26] ), .Z(n4941) );
  CIVX2 U4076 ( .A(\reg_mem[29][26] ), .Z(n4971) );
  CMXI2X1 U4077 ( .A0(n4941), .A1(n4971), .S(n2104), .Z(n2636) );
  CIVX2 U4078 ( .A(\reg_mem[15][26] ), .Z(n4943) );
  CIVX2 U4079 ( .A(\reg_mem[31][26] ), .Z(n4973) );
  CMXI2X1 U4080 ( .A0(n4943), .A1(n4973), .S(n2087), .Z(n2635) );
  CMXI2X1 U4081 ( .A0(n2636), .A1(n2635), .S(n2189), .Z(n2637) );
  CIVX2 U4082 ( .A(\reg_mem[0][26] ), .Z(n4922) );
  CIVX2 U4083 ( .A(\reg_mem[16][26] ), .Z(n4952) );
  CMXI2X1 U4084 ( .A0(n4922), .A1(n4952), .S(n2091), .Z(n2641) );
  CIVX2 U4085 ( .A(\reg_mem[2][26] ), .Z(n4924) );
  CIVX2 U4086 ( .A(\reg_mem[18][26] ), .Z(n4954) );
  CMXI2X1 U4087 ( .A0(n4924), .A1(n4954), .S(n2080), .Z(n2640) );
  CIVX2 U4088 ( .A(\reg_mem[4][26] ), .Z(n4928) );
  CIVX2 U4089 ( .A(\reg_mem[20][26] ), .Z(n4958) );
  CMXI2X1 U4090 ( .A0(n4928), .A1(n4958), .S(n2080), .Z(n2643) );
  CIVX2 U4091 ( .A(\reg_mem[6][26] ), .Z(n4930) );
  CIVX2 U4092 ( .A(\reg_mem[22][26] ), .Z(n4960) );
  CMXI2X1 U4093 ( .A0(n4930), .A1(n4960), .S(n2097), .Z(n2642) );
  CIVX2 U4094 ( .A(n3631), .Z(n2694) );
  CIVX2 U4095 ( .A(\reg_mem[1][26] ), .Z(n4921) );
  CIVX2 U4096 ( .A(\reg_mem[17][26] ), .Z(n4951) );
  CMXI2X1 U4097 ( .A0(n4921), .A1(n4951), .S(n2081), .Z(n2648) );
  CIVX2 U4098 ( .A(\reg_mem[3][26] ), .Z(n4923) );
  CIVX2 U4099 ( .A(\reg_mem[19][26] ), .Z(n4953) );
  CMXI2X1 U4100 ( .A0(n4923), .A1(n4953), .S(n2092), .Z(n2647) );
  CMXI2X1 U4101 ( .A0(n2648), .A1(n2647), .S(n2178), .Z(n2652) );
  CIVX2 U4102 ( .A(\reg_mem[5][26] ), .Z(n4927) );
  CIVX2 U4103 ( .A(\reg_mem[21][26] ), .Z(n4957) );
  CMXI2X1 U4104 ( .A0(n4927), .A1(n4957), .S(n2090), .Z(n2650) );
  CIVX2 U4105 ( .A(\reg_mem[7][26] ), .Z(n4929) );
  CIVX2 U4106 ( .A(\reg_mem[23][26] ), .Z(n4959) );
  CMXI2X1 U4107 ( .A0(n4929), .A1(n4959), .S(n2096), .Z(n2649) );
  CMXI2X1 U4108 ( .A0(n2650), .A1(n2649), .S(n2180), .Z(n2651) );
  CMXI2X1 U4109 ( .A0(n2652), .A1(n2651), .S(net87266), .Z(n2653) );
  CIVX2 U4110 ( .A(n3623), .Z(n2702) );
  CIVX2 U4111 ( .A(\reg_mem[8][26] ), .Z(n4936) );
  CIVX2 U4112 ( .A(\reg_mem[24][26] ), .Z(n4966) );
  CIVX2 U4113 ( .A(\reg_mem[10][26] ), .Z(n4938) );
  CIVX2 U4114 ( .A(\reg_mem[26][26] ), .Z(n4968) );
  CIVX2 U4115 ( .A(\reg_mem[12][26] ), .Z(n4942) );
  CIVX2 U4116 ( .A(\reg_mem[28][26] ), .Z(n4972) );
  CIVX2 U4117 ( .A(\reg_mem[14][26] ), .Z(n4944) );
  CIVX2 U4118 ( .A(\reg_mem[30][26] ), .Z(n4974) );
  CMXI2X1 U4119 ( .A0(n4944), .A1(n4974), .S(n2083), .Z(n2656) );
  CIVX2 U4120 ( .A(N121), .Z(n2671) );
  CIVX2 U4121 ( .A(\reg_mem[9][25] ), .Z(n4873) );
  CIVX2 U4122 ( .A(\reg_mem[25][25] ), .Z(n4903) );
  CMXI2X1 U4123 ( .A0(n4873), .A1(n4903), .S(n2089), .Z(n2673) );
  CIVX2 U4124 ( .A(\reg_mem[11][25] ), .Z(n4875) );
  CIVX2 U4125 ( .A(\reg_mem[27][25] ), .Z(n4905) );
  CMXI2X1 U4126 ( .A0(n4875), .A1(n4905), .S(n2088), .Z(n2672) );
  CMXI2X1 U4127 ( .A0(n2673), .A1(n2672), .S(n2177), .Z(n2677) );
  CIVX2 U4128 ( .A(\reg_mem[13][25] ), .Z(n4879) );
  CIVX2 U4129 ( .A(\reg_mem[29][25] ), .Z(n4909) );
  CMXI2X1 U4130 ( .A0(n4879), .A1(n4909), .S(n2098), .Z(n2675) );
  CIVX2 U4131 ( .A(\reg_mem[15][25] ), .Z(n4881) );
  CIVX2 U4132 ( .A(\reg_mem[31][25] ), .Z(n4911) );
  CIVX2 U4133 ( .A(\reg_mem[0][25] ), .Z(n4860) );
  CIVX2 U4134 ( .A(\reg_mem[16][25] ), .Z(n4890) );
  CIVX2 U4135 ( .A(\reg_mem[2][25] ), .Z(n4862) );
  CIVX2 U4136 ( .A(\reg_mem[18][25] ), .Z(n4892) );
  CIVX2 U4137 ( .A(\reg_mem[4][25] ), .Z(n4866) );
  CIVX2 U4138 ( .A(\reg_mem[20][25] ), .Z(n4896) );
  CMXI2X1 U4139 ( .A0(n4866), .A1(n4896), .S(n2090), .Z(n2682) );
  CIVX2 U4140 ( .A(\reg_mem[6][25] ), .Z(n4868) );
  CIVX2 U4141 ( .A(\reg_mem[22][25] ), .Z(n4898) );
  CMXI2X1 U4142 ( .A0(n4868), .A1(n4898), .S(n2090), .Z(n2681) );
  CIVX2 U4143 ( .A(\reg_mem[1][25] ), .Z(n4859) );
  CIVX2 U4144 ( .A(\reg_mem[17][25] ), .Z(n4889) );
  CMXI2X1 U4145 ( .A0(n4859), .A1(n4889), .S(n2099), .Z(n2688) );
  CIVX2 U4146 ( .A(\reg_mem[3][25] ), .Z(n4861) );
  CIVX2 U4147 ( .A(\reg_mem[19][25] ), .Z(n4891) );
  CIVX2 U4148 ( .A(\reg_mem[5][25] ), .Z(n4865) );
  CIVX2 U4149 ( .A(\reg_mem[21][25] ), .Z(n4895) );
  CMXI2X1 U4150 ( .A0(n4865), .A1(n4895), .S(n2085), .Z(n2690) );
  CIVX2 U4151 ( .A(\reg_mem[7][25] ), .Z(n4867) );
  CIVX2 U4152 ( .A(\reg_mem[23][25] ), .Z(n4897) );
  CMXI2X1 U4153 ( .A0(n4867), .A1(n4897), .S(n2091), .Z(n2689) );
  CMXI2X1 U4154 ( .A0(n2690), .A1(n2689), .S(n2185), .Z(n2691) );
  CMXI2X1 U4155 ( .A0(n2692), .A1(n2691), .S(net87262), .Z(n2693) );
  CIVX2 U4156 ( .A(\reg_mem[8][25] ), .Z(n4874) );
  CIVX2 U4157 ( .A(\reg_mem[24][25] ), .Z(n4904) );
  CIVX2 U4158 ( .A(\reg_mem[10][25] ), .Z(n4876) );
  CIVX2 U4159 ( .A(\reg_mem[26][25] ), .Z(n4906) );
  CMXI2X1 U4160 ( .A0(n4876), .A1(n4906), .S(n2084), .Z(n2695) );
  CMXI2X1 U4161 ( .A0(n2696), .A1(n2695), .S(n2181), .Z(n2700) );
  CIVX2 U4162 ( .A(\reg_mem[12][25] ), .Z(n4880) );
  CIVX2 U4163 ( .A(\reg_mem[28][25] ), .Z(n4910) );
  CMXI2X1 U4164 ( .A0(n4880), .A1(n4910), .S(n2085), .Z(n2698) );
  CIVX2 U4165 ( .A(\reg_mem[14][25] ), .Z(n4882) );
  CIVX2 U4166 ( .A(\reg_mem[30][25] ), .Z(n4912) );
  CMXI2X1 U4167 ( .A0(n4882), .A1(n4912), .S(n2083), .Z(n2697) );
  CND2IX1 U4168 ( .B(n2711), .A(n2710), .Z(alu_op_c[25]) );
  CIVX2 U4169 ( .A(n2712), .Z(n2715) );
  CND2IX1 U4170 ( .B(n3181), .A(N161), .Z(n2713) );
  CMXI2X1 U4171 ( .A0(\reg_mem[0][24] ), .A1(\reg_mem[16][24] ), .S(n2082), 
        .Z(n2719) );
  CMXI2X1 U4172 ( .A0(\reg_mem[2][24] ), .A1(\reg_mem[18][24] ), .S(n2083), 
        .Z(n2718) );
  CMXI2X1 U4173 ( .A0(n2719), .A1(n2718), .S(n2176), .Z(n2723) );
  CMXI2X1 U4174 ( .A0(\reg_mem[4][24] ), .A1(\reg_mem[20][24] ), .S(n2084), 
        .Z(n2721) );
  CMXI2X1 U4175 ( .A0(\reg_mem[6][24] ), .A1(\reg_mem[22][24] ), .S(n2089), 
        .Z(n2720) );
  CMXI2X1 U4176 ( .A0(n2723), .A1(n2722), .S(net87278), .Z(n2731) );
  CMXI2X1 U4177 ( .A0(\reg_mem[8][24] ), .A1(\reg_mem[24][24] ), .S(n2081), 
        .Z(n2725) );
  CMXI2X1 U4178 ( .A0(\reg_mem[10][24] ), .A1(\reg_mem[26][24] ), .S(n2091), 
        .Z(n2724) );
  CMXI2X1 U4179 ( .A0(\reg_mem[12][24] ), .A1(\reg_mem[28][24] ), .S(n2081), 
        .Z(n2727) );
  CMXI2X1 U4180 ( .A0(\reg_mem[14][24] ), .A1(\reg_mem[30][24] ), .S(n2102), 
        .Z(n2726) );
  CMXI2X1 U4181 ( .A0(n2729), .A1(n2728), .S(net87279), .Z(n2730) );
  CMXI2X1 U4182 ( .A0(\reg_mem[1][24] ), .A1(\reg_mem[17][24] ), .S(n2080), 
        .Z(n2733) );
  CMXI2X1 U4183 ( .A0(\reg_mem[5][24] ), .A1(\reg_mem[21][24] ), .S(n2080), 
        .Z(n2735) );
  CMXI2X1 U4184 ( .A0(\reg_mem[7][24] ), .A1(\reg_mem[23][24] ), .S(n2080), 
        .Z(n2734) );
  CMXI2X1 U4185 ( .A0(\reg_mem[9][24] ), .A1(\reg_mem[25][24] ), .S(n2103), 
        .Z(n2739) );
  CMXI2X1 U4186 ( .A0(\reg_mem[11][24] ), .A1(\reg_mem[27][24] ), .S(n2105), 
        .Z(n2738) );
  CMXI2X1 U4187 ( .A0(\reg_mem[13][24] ), .A1(\reg_mem[29][24] ), .S(n2105), 
        .Z(n2741) );
  CMXI2X1 U4188 ( .A0(\reg_mem[15][24] ), .A1(\reg_mem[31][24] ), .S(n2081), 
        .Z(n2740) );
  CMXI2X1 U4189 ( .A0(n2741), .A1(n2740), .S(n2189), .Z(n2742) );
  CMXI2X1 U4190 ( .A0(n2743), .A1(n2742), .S(net87247), .Z(n2744) );
  CMXI2X1 U4191 ( .A0(\reg_mem[0][23] ), .A1(\reg_mem[8][23] ), .S(net87538), 
        .Z(n2749) );
  CMXI2X1 U4192 ( .A0(\reg_mem[2][23] ), .A1(\reg_mem[10][23] ), .S(net87533), 
        .Z(n2748) );
  CMXI2X1 U4193 ( .A0(n2749), .A1(n2748), .S(n2191), .Z(n2753) );
  CMXI2X1 U4194 ( .A0(\reg_mem[4][23] ), .A1(\reg_mem[12][23] ), .S(net87529), 
        .Z(n2751) );
  CMXI2X1 U4195 ( .A0(\reg_mem[6][23] ), .A1(\reg_mem[14][23] ), .S(net87520), 
        .Z(n2750) );
  CMXI2X1 U4196 ( .A0(n2751), .A1(n2750), .S(n2193), .Z(n2752) );
  CMXI2X1 U4197 ( .A0(n2753), .A1(n2752), .S(net87278), .Z(n2761) );
  CMXI2X1 U4198 ( .A0(\reg_mem[1][23] ), .A1(\reg_mem[9][23] ), .S(net87544), 
        .Z(n2755) );
  CMXI2X1 U4199 ( .A0(\reg_mem[3][23] ), .A1(\reg_mem[11][23] ), .S(net87540), 
        .Z(n2754) );
  CMXI2X1 U4200 ( .A0(n2755), .A1(n2754), .S(n2197), .Z(n2759) );
  CMXI2X1 U4201 ( .A0(\reg_mem[5][23] ), .A1(\reg_mem[13][23] ), .S(net87523), 
        .Z(n2757) );
  CMXI2X1 U4202 ( .A0(n2757), .A1(n2756), .S(n2199), .Z(n2758) );
  CMXI2X1 U4203 ( .A0(n2759), .A1(n2758), .S(net87278), .Z(n2760) );
  CMXI2X1 U4204 ( .A0(n2761), .A1(n2760), .S(net87395), .Z(n2777) );
  CMXI2X1 U4205 ( .A0(\reg_mem[16][23] ), .A1(\reg_mem[24][23] ), .S(net87520), 
        .Z(n2763) );
  CMXI2X1 U4206 ( .A0(\reg_mem[18][23] ), .A1(\reg_mem[26][23] ), .S(net87540), 
        .Z(n2762) );
  CMXI2X1 U4207 ( .A0(n2763), .A1(n2762), .S(n2194), .Z(n2767) );
  CMXI2X1 U4208 ( .A0(\reg_mem[20][23] ), .A1(\reg_mem[28][23] ), .S(net87530), 
        .Z(n2765) );
  CMXI2X1 U4209 ( .A0(\reg_mem[22][23] ), .A1(\reg_mem[30][23] ), .S(net87522), 
        .Z(n2764) );
  CMXI2X1 U4210 ( .A0(n2765), .A1(n2764), .S(n2195), .Z(n2766) );
  CMXI2X1 U4211 ( .A0(n2767), .A1(n2766), .S(net87268), .Z(n2775) );
  CMXI2X1 U4212 ( .A0(\reg_mem[17][23] ), .A1(\reg_mem[25][23] ), .S(net87533), 
        .Z(n2769) );
  CMXI2X1 U4213 ( .A0(\reg_mem[19][23] ), .A1(\reg_mem[27][23] ), .S(net87525), 
        .Z(n2768) );
  CMXI2X1 U4214 ( .A0(n2769), .A1(n2768), .S(n2183), .Z(n2773) );
  CMXI2X1 U4215 ( .A0(\reg_mem[21][23] ), .A1(\reg_mem[29][23] ), .S(net87519), 
        .Z(n2771) );
  CMXI2X1 U4216 ( .A0(\reg_mem[23][23] ), .A1(\reg_mem[31][23] ), .S(net87526), 
        .Z(n2770) );
  CMXI2X1 U4217 ( .A0(n2771), .A1(n2770), .S(n2185), .Z(n2772) );
  CMXI2X1 U4218 ( .A0(n2773), .A1(n2772), .S(net87273), .Z(n2774) );
  CMXI2X1 U4219 ( .A0(n2775), .A1(n2774), .S(net87397), .Z(n2776) );
  CMXI2X1 U4220 ( .A0(n2777), .A1(n2776), .S(n2088), .Z(n2778) );
  CIVX2 U4221 ( .A(n2779), .Z(n2782) );
  CND2IX1 U4222 ( .B(n3181), .A(N160), .Z(n2780) );
  CND2IX1 U4223 ( .B(n3181), .A(N159), .Z(n2788) );
  CIVX2 U4224 ( .A(\reg_mem[17][22] ), .Z(n4739) );
  CIVX2 U4225 ( .A(\reg_mem[25][22] ), .Z(n4753) );
  CMXI2X1 U4226 ( .A0(n4739), .A1(n4753), .S(net87522), .Z(n2791) );
  CIVX2 U4227 ( .A(\reg_mem[19][22] ), .Z(n4741) );
  CIVX2 U4228 ( .A(\reg_mem[27][22] ), .Z(n4755) );
  CMXI2X1 U4229 ( .A0(n4741), .A1(n4755), .S(net87525), .Z(n2790) );
  CMXI2X1 U4230 ( .A0(n2791), .A1(n2790), .S(n2184), .Z(n2795) );
  CIVX2 U4231 ( .A(\reg_mem[21][22] ), .Z(n4745) );
  CIVX2 U4232 ( .A(\reg_mem[29][22] ), .Z(n4759) );
  CMXI2X1 U4233 ( .A0(n4745), .A1(n4759), .S(net87544), .Z(n2793) );
  CIVX2 U4234 ( .A(\reg_mem[23][22] ), .Z(n4747) );
  CIVX2 U4235 ( .A(\reg_mem[31][22] ), .Z(n4761) );
  CMXI2X1 U4236 ( .A0(n4747), .A1(n4761), .S(net87526), .Z(n2792) );
  CMXI2X1 U4237 ( .A0(n2793), .A1(n2792), .S(n2180), .Z(n2794) );
  CIVX2 U4238 ( .A(\reg_mem[0][22] ), .Z(n4710) );
  CIVX2 U4239 ( .A(\reg_mem[8][22] ), .Z(n4724) );
  CMXI2X1 U4240 ( .A0(n4710), .A1(n4724), .S(net87541), .Z(n2799) );
  CIVX2 U4241 ( .A(\reg_mem[2][22] ), .Z(n4712) );
  CIVX2 U4242 ( .A(\reg_mem[10][22] ), .Z(n4726) );
  CMXI2X1 U4243 ( .A0(n4712), .A1(n4726), .S(net87532), .Z(n2798) );
  CMXI2X1 U4244 ( .A0(n2799), .A1(n2798), .S(n2178), .Z(n2803) );
  CIVX2 U4245 ( .A(\reg_mem[4][22] ), .Z(n4716) );
  CIVX2 U4246 ( .A(\reg_mem[12][22] ), .Z(n4730) );
  CMXI2X1 U4247 ( .A0(n4716), .A1(n4730), .S(net87519), .Z(n2801) );
  CIVX2 U4248 ( .A(\reg_mem[6][22] ), .Z(n4718) );
  CIVX2 U4249 ( .A(\reg_mem[14][22] ), .Z(n4732) );
  CMXI2X1 U4250 ( .A0(n2803), .A1(n2802), .S(net87247), .Z(n2804) );
  CIVX2 U4251 ( .A(\reg_mem[16][22] ), .Z(n4740) );
  CIVX2 U4252 ( .A(\reg_mem[24][22] ), .Z(n4754) );
  CMXI2X1 U4253 ( .A0(n4740), .A1(n4754), .S(net87522), .Z(n2807) );
  CIVX2 U4254 ( .A(\reg_mem[18][22] ), .Z(n4742) );
  CIVX2 U4255 ( .A(\reg_mem[26][22] ), .Z(n4756) );
  CMXI2X1 U4256 ( .A0(n4742), .A1(n4756), .S(net87520), .Z(n2806) );
  CMXI2X1 U4257 ( .A0(n2807), .A1(n2806), .S(n2166), .Z(n2811) );
  CIVX2 U4258 ( .A(\reg_mem[20][22] ), .Z(n4746) );
  CIVX2 U4259 ( .A(\reg_mem[28][22] ), .Z(n4760) );
  CMXI2X1 U4260 ( .A0(n4746), .A1(n4760), .S(net87519), .Z(n2809) );
  CIVX2 U4261 ( .A(\reg_mem[22][22] ), .Z(n4748) );
  CIVX2 U4262 ( .A(\reg_mem[30][22] ), .Z(n4762) );
  CMXI2X1 U4263 ( .A0(n4748), .A1(n4762), .S(net87542), .Z(n2808) );
  CMXI2X1 U4264 ( .A0(n2809), .A1(n2808), .S(n2182), .Z(n2810) );
  CMXI2X1 U4265 ( .A0(n2811), .A1(n2810), .S(net87276), .Z(n2812) );
  CIVX2 U4266 ( .A(\reg_mem[1][22] ), .Z(n4709) );
  CIVX2 U4267 ( .A(\reg_mem[9][22] ), .Z(n4723) );
  CIVX2 U4268 ( .A(\reg_mem[3][22] ), .Z(n4711) );
  CIVX2 U4269 ( .A(\reg_mem[11][22] ), .Z(n4725) );
  CMXI2X1 U4270 ( .A0(n4711), .A1(n4725), .S(net87521), .Z(n2814) );
  CIVX2 U4271 ( .A(\reg_mem[5][22] ), .Z(n4715) );
  CIVX2 U4272 ( .A(\reg_mem[13][22] ), .Z(n4729) );
  CMXI2X1 U4273 ( .A0(n4715), .A1(n4729), .S(net87540), .Z(n2817) );
  CIVX2 U4274 ( .A(\reg_mem[7][22] ), .Z(n4717) );
  CIVX2 U4275 ( .A(\reg_mem[15][22] ), .Z(n4731) );
  CMXI2X1 U4276 ( .A0(n4717), .A1(n4731), .S(net87540), .Z(n2816) );
  CND2IX1 U4277 ( .B(n2828), .A(n2827), .Z(n5245) );
  CIVX2 U4278 ( .A(\reg_mem[5][21] ), .Z(n4653) );
  CIVX2 U4279 ( .A(\reg_mem[21][21] ), .Z(n4683) );
  CMXI2X1 U4280 ( .A0(n4653), .A1(n4683), .S(n2102), .Z(n2833) );
  CIVX2 U4281 ( .A(\reg_mem[7][21] ), .Z(n4655) );
  CIVX2 U4282 ( .A(\reg_mem[23][21] ), .Z(n4685) );
  CND2IX1 U4283 ( .B(n3649), .A(n2834), .Z(n2843) );
  CIVX2 U4284 ( .A(\reg_mem[9][21] ), .Z(n4661) );
  CIVX2 U4285 ( .A(\reg_mem[25][21] ), .Z(n4691) );
  CMXI2X1 U4286 ( .A0(n4661), .A1(n4691), .S(n2085), .Z(n2836) );
  CIVX2 U4287 ( .A(\reg_mem[11][21] ), .Z(n4663) );
  CIVX2 U4288 ( .A(\reg_mem[27][21] ), .Z(n4693) );
  CIVX2 U4289 ( .A(\reg_mem[13][21] ), .Z(n4667) );
  CIVX2 U4290 ( .A(\reg_mem[29][21] ), .Z(n4697) );
  CIVX2 U4291 ( .A(\reg_mem[15][21] ), .Z(n4669) );
  CIVX2 U4292 ( .A(\reg_mem[31][21] ), .Z(n4699) );
  CMXI2X1 U4293 ( .A0(n2839), .A1(n2838), .S(n2166), .Z(n2840) );
  CIVX2 U4294 ( .A(\reg_mem[8][21] ), .Z(n4662) );
  CIVX2 U4295 ( .A(\reg_mem[24][21] ), .Z(n4692) );
  CMXI2X1 U4296 ( .A0(n4662), .A1(n4692), .S(n2082), .Z(n2845) );
  CIVX2 U4297 ( .A(\reg_mem[10][21] ), .Z(n4664) );
  CIVX2 U4298 ( .A(\reg_mem[26][21] ), .Z(n4694) );
  CIVX2 U4299 ( .A(\reg_mem[12][21] ), .Z(n4668) );
  CIVX2 U4300 ( .A(\reg_mem[28][21] ), .Z(n4698) );
  CMXI2X1 U4301 ( .A0(n4668), .A1(n4698), .S(n2091), .Z(n2848) );
  CIVX2 U4302 ( .A(\reg_mem[14][21] ), .Z(n4670) );
  CIVX2 U4303 ( .A(\reg_mem[30][21] ), .Z(n4700) );
  CMXI2X1 U4304 ( .A0(n4670), .A1(n4700), .S(n2100), .Z(n2847) );
  CMXI2X1 U4305 ( .A0(n2848), .A1(n2847), .S(n1469), .Z(n2849) );
  CND2IX1 U4306 ( .B(n3667), .A(n2849), .Z(n2854) );
  CIVX2 U4307 ( .A(\reg_mem[1][21] ), .Z(n4647) );
  CIVX2 U4308 ( .A(\reg_mem[17][21] ), .Z(n4677) );
  CMXI2X1 U4309 ( .A0(n4647), .A1(n4677), .S(n2092), .Z(n2851) );
  CIVX2 U4310 ( .A(\reg_mem[3][21] ), .Z(n4649) );
  CIVX2 U4311 ( .A(\reg_mem[19][21] ), .Z(n4679) );
  CMXI2X1 U4312 ( .A0(n4649), .A1(n4679), .S(n2105), .Z(n2850) );
  CMXI2X1 U4313 ( .A0(n2851), .A1(n2850), .S(n2193), .Z(n2852) );
  CND2IX1 U4314 ( .B(n3671), .A(n2852), .Z(n2853) );
  CMXI2X1 U4315 ( .A0(\reg_mem[0][21] ), .A1(\reg_mem[16][21] ), .S(n2091), 
        .Z(n2857) );
  CMXI2X1 U4316 ( .A0(\reg_mem[2][21] ), .A1(\reg_mem[18][21] ), .S(n2022), 
        .Z(n2856) );
  CMXI2X1 U4317 ( .A0(n2857), .A1(n2856), .S(n1469), .Z(n2861) );
  CMXI2X1 U4318 ( .A0(n2859), .A1(n2858), .S(n2180), .Z(n2860) );
  CMXI2X1 U4319 ( .A0(\reg_mem[0][20] ), .A1(\reg_mem[8][20] ), .S(net87530), 
        .Z(n2871) );
  CMXI2X1 U4320 ( .A0(\reg_mem[2][20] ), .A1(\reg_mem[10][20] ), .S(net87541), 
        .Z(n2870) );
  CMXI2X1 U4321 ( .A0(n2871), .A1(n2870), .S(n2190), .Z(n2875) );
  CMXI2X1 U4322 ( .A0(\reg_mem[4][20] ), .A1(\reg_mem[12][20] ), .S(net87542), 
        .Z(n2873) );
  CMXI2X1 U4323 ( .A0(\reg_mem[6][20] ), .A1(\reg_mem[14][20] ), .S(net87531), 
        .Z(n2872) );
  CMXI2X1 U4324 ( .A0(n2873), .A1(n2872), .S(n2192), .Z(n2874) );
  CMXI2X1 U4325 ( .A0(n2875), .A1(n2874), .S(net87281), .Z(n2883) );
  CMXI2X1 U4326 ( .A0(\reg_mem[1][20] ), .A1(\reg_mem[9][20] ), .S(net87532), 
        .Z(n2877) );
  CMXI2X1 U4327 ( .A0(\reg_mem[3][20] ), .A1(\reg_mem[11][20] ), .S(net87529), 
        .Z(n2876) );
  CMXI2X1 U4328 ( .A0(n2877), .A1(n2876), .S(n2196), .Z(n2881) );
  CMXI2X1 U4329 ( .A0(\reg_mem[7][20] ), .A1(\reg_mem[15][20] ), .S(net87521), 
        .Z(n2878) );
  CMXI2X1 U4330 ( .A0(n2881), .A1(n2880), .S(n1480), .Z(n2882) );
  CMXI2X1 U4331 ( .A0(n2883), .A1(n2882), .S(net87394), .Z(n2898) );
  CMXI2X1 U4332 ( .A0(\reg_mem[18][20] ), .A1(\reg_mem[26][20] ), .S(net87531), 
        .Z(n2884) );
  CMXI2X1 U4333 ( .A0(n2885), .A1(n2884), .S(n2162), .Z(n2888) );
  CMXI2X1 U4334 ( .A0(\reg_mem[21][20] ), .A1(\reg_mem[29][20] ), .S(net87522), 
        .Z(n2892) );
  CMXI2X1 U4335 ( .A0(\reg_mem[23][20] ), .A1(\reg_mem[31][20] ), .S(net87522), 
        .Z(n2891) );
  CMXI2X1 U4336 ( .A0(n2892), .A1(n2891), .S(n2184), .Z(n2893) );
  CMXI2X1 U4337 ( .A0(n2894), .A1(n2893), .S(net87247), .Z(n2895) );
  CMXI2X1 U4338 ( .A0(n2898), .A1(n2897), .S(n2022), .Z(n2899) );
  CIVX2 U4339 ( .A(N116), .Z(n2902) );
  COND3X1 U4340 ( .A(n2123), .B(n2902), .C(n2901), .D(n2900), .Z(n2906) );
  CND2IX1 U4341 ( .B(n2904), .A(n2903), .Z(N289) );
  CND2IX1 U4342 ( .B(n2906), .A(n2905), .Z(alu_op_c[20]) );
  CMXI2X1 U4343 ( .A0(\reg_mem[0][19] ), .A1(\reg_mem[8][19] ), .S(net87520), 
        .Z(n2911) );
  CMXI2X1 U4344 ( .A0(\reg_mem[4][19] ), .A1(\reg_mem[12][19] ), .S(net87542), 
        .Z(n2913) );
  CMXI2X1 U4345 ( .A0(\reg_mem[6][19] ), .A1(\reg_mem[14][19] ), .S(net87542), 
        .Z(n2912) );
  CMXI2X1 U4346 ( .A0(n2913), .A1(n2912), .S(n2185), .Z(n2914) );
  CMXI2X1 U4347 ( .A0(n2915), .A1(n2914), .S(net87278), .Z(n2923) );
  CMXI2X1 U4348 ( .A0(\reg_mem[1][19] ), .A1(\reg_mem[9][19] ), .S(net87520), 
        .Z(n2917) );
  CMXI2X1 U4349 ( .A0(\reg_mem[3][19] ), .A1(\reg_mem[11][19] ), .S(net87530), 
        .Z(n2916) );
  CMXI2X1 U4350 ( .A0(n2917), .A1(n2916), .S(n1469), .Z(n2921) );
  CMXI2X1 U4351 ( .A0(\reg_mem[5][19] ), .A1(\reg_mem[13][19] ), .S(net87538), 
        .Z(n2919) );
  CMXI2X1 U4352 ( .A0(\reg_mem[7][19] ), .A1(\reg_mem[15][19] ), .S(net87531), 
        .Z(n2918) );
  CMXI2X1 U4353 ( .A0(n2919), .A1(n2918), .S(n2177), .Z(n2920) );
  CMXI2X1 U4354 ( .A0(n2921), .A1(n2920), .S(net87269), .Z(n2922) );
  CMXI2X1 U4355 ( .A0(\reg_mem[16][19] ), .A1(\reg_mem[24][19] ), .S(net87531), 
        .Z(n2925) );
  CMXI2X1 U4356 ( .A0(\reg_mem[18][19] ), .A1(\reg_mem[26][19] ), .S(net87524), 
        .Z(n2924) );
  CMXI2X1 U4357 ( .A0(n2925), .A1(n2924), .S(n2197), .Z(n2929) );
  CMXI2X1 U4358 ( .A0(\reg_mem[20][19] ), .A1(\reg_mem[28][19] ), .S(net87533), 
        .Z(n2927) );
  CMXI2X1 U4359 ( .A0(\reg_mem[22][19] ), .A1(\reg_mem[30][19] ), .S(net87541), 
        .Z(n2926) );
  CMXI2X1 U4360 ( .A0(n2927), .A1(n2926), .S(n2192), .Z(n2928) );
  CMXI2X1 U4361 ( .A0(n2929), .A1(n2928), .S(net87261), .Z(n2937) );
  CMXI2X1 U4362 ( .A0(\reg_mem[17][19] ), .A1(\reg_mem[25][19] ), .S(net87529), 
        .Z(n2931) );
  CMXI2X1 U4363 ( .A0(\reg_mem[19][19] ), .A1(\reg_mem[27][19] ), .S(net87532), 
        .Z(n2930) );
  CMXI2X1 U4364 ( .A0(n2931), .A1(n2930), .S(n2183), .Z(n2935) );
  CMXI2X1 U4365 ( .A0(\reg_mem[21][19] ), .A1(\reg_mem[29][19] ), .S(net87541), 
        .Z(n2933) );
  CMXI2X1 U4366 ( .A0(\reg_mem[23][19] ), .A1(\reg_mem[31][19] ), .S(net87540), 
        .Z(n2932) );
  CMXI2X1 U4367 ( .A0(n2935), .A1(n2934), .S(n1391), .Z(n2936) );
  CMXI2X1 U4368 ( .A0(n2937), .A1(n2936), .S(net87402), .Z(n2938) );
  CMXI2X1 U4369 ( .A0(n2939), .A1(n2938), .S(n2094), .Z(n2941) );
  CMXI2X1 U4370 ( .A0(n2941), .A1(n2940), .S(n1533), .Z(N288) );
  CANR2X1 U4371 ( .A(N187), .B(n3704), .C(N155), .D(n3701), .Z(n2944) );
  CMXI2X1 U4372 ( .A0(\reg_mem[0][18] ), .A1(\reg_mem[16][18] ), .S(n2097), 
        .Z(n2946) );
  CMXI2X1 U4373 ( .A0(\reg_mem[2][18] ), .A1(\reg_mem[18][18] ), .S(n2100), 
        .Z(n2945) );
  CMXI2X1 U4374 ( .A0(n2946), .A1(n2945), .S(n2199), .Z(n2950) );
  CMXI2X1 U4375 ( .A0(\reg_mem[6][18] ), .A1(\reg_mem[22][18] ), .S(n2084), 
        .Z(n2947) );
  CMXI2X1 U4376 ( .A0(n2950), .A1(n2949), .S(net87248), .Z(n2958) );
  CMXI2X1 U4377 ( .A0(\reg_mem[8][18] ), .A1(\reg_mem[24][18] ), .S(n2091), 
        .Z(n2952) );
  CMXI2X1 U4378 ( .A0(\reg_mem[10][18] ), .A1(\reg_mem[26][18] ), .S(n2104), 
        .Z(n2951) );
  CMXI2X1 U4379 ( .A0(n2952), .A1(n2951), .S(n2179), .Z(n2956) );
  CMXI2X1 U4380 ( .A0(\reg_mem[12][18] ), .A1(\reg_mem[28][18] ), .S(n2087), 
        .Z(n2954) );
  CMXI2X1 U4381 ( .A0(\reg_mem[14][18] ), .A1(\reg_mem[30][18] ), .S(n2100), 
        .Z(n2953) );
  CMXI2X1 U4382 ( .A0(n2954), .A1(n2953), .S(n2162), .Z(n2955) );
  CMXI2X1 U4383 ( .A0(\reg_mem[1][18] ), .A1(\reg_mem[17][18] ), .S(n2092), 
        .Z(n2960) );
  CMXI2X1 U4384 ( .A0(\reg_mem[3][18] ), .A1(\reg_mem[19][18] ), .S(n2083), 
        .Z(n2959) );
  CMXI2X1 U4385 ( .A0(n2960), .A1(n2959), .S(n2196), .Z(n2964) );
  CMXI2X1 U4386 ( .A0(\reg_mem[5][18] ), .A1(\reg_mem[21][18] ), .S(n2096), 
        .Z(n2962) );
  CMXI2X1 U4387 ( .A0(\reg_mem[7][18] ), .A1(\reg_mem[23][18] ), .S(n2104), 
        .Z(n2961) );
  CMXI2X1 U4388 ( .A0(n2964), .A1(n2963), .S(n1385), .Z(n2972) );
  CMXI2X1 U4389 ( .A0(\reg_mem[9][18] ), .A1(\reg_mem[25][18] ), .S(n2099), 
        .Z(n2966) );
  CMXI2X1 U4390 ( .A0(\reg_mem[11][18] ), .A1(\reg_mem[27][18] ), .S(n2101), 
        .Z(n2965) );
  CMXI2X1 U4391 ( .A0(\reg_mem[13][18] ), .A1(\reg_mem[29][18] ), .S(n2095), 
        .Z(n2968) );
  CIVX2 U4392 ( .A(N113), .Z(n2974) );
  CIVX2 U4393 ( .A(N81), .Z(n2973) );
  CANR2X1 U4394 ( .A(N186), .B(n3704), .C(N154), .D(n3701), .Z(n2975) );
  CND2IX1 U4395 ( .B(n2976), .A(n2975), .Z(alu_op_c[17]) );
  CMXI2X1 U4396 ( .A0(\reg_mem[0][17] ), .A1(\reg_mem[8][17] ), .S(net87542), 
        .Z(n2978) );
  CMXI2X1 U4397 ( .A0(\reg_mem[2][17] ), .A1(\reg_mem[10][17] ), .S(net87530), 
        .Z(n2977) );
  CMXI2X1 U4398 ( .A0(n2978), .A1(n2977), .S(n2198), .Z(n2982) );
  CMXI2X1 U4399 ( .A0(\reg_mem[4][17] ), .A1(\reg_mem[12][17] ), .S(net87541), 
        .Z(n2980) );
  CMXI2X1 U4400 ( .A0(\reg_mem[6][17] ), .A1(\reg_mem[14][17] ), .S(net87541), 
        .Z(n2979) );
  CMXI2X1 U4401 ( .A0(n2982), .A1(n2981), .S(n1385), .Z(n2990) );
  CMXI2X1 U4402 ( .A0(\reg_mem[1][17] ), .A1(\reg_mem[9][17] ), .S(net87521), 
        .Z(n2984) );
  CMXI2X1 U4403 ( .A0(\reg_mem[3][17] ), .A1(\reg_mem[11][17] ), .S(net87545), 
        .Z(n2983) );
  CMXI2X1 U4404 ( .A0(n2984), .A1(n2983), .S(n2178), .Z(n2988) );
  CMXI2X1 U4405 ( .A0(\reg_mem[5][17] ), .A1(\reg_mem[13][17] ), .S(net87538), 
        .Z(n2986) );
  CMXI2X1 U4406 ( .A0(\reg_mem[7][17] ), .A1(\reg_mem[15][17] ), .S(net87545), 
        .Z(n2985) );
  CMXI2X1 U4407 ( .A0(\reg_mem[16][17] ), .A1(\reg_mem[24][17] ), .S(net87545), 
        .Z(n2992) );
  CMXI2X1 U4408 ( .A0(\reg_mem[18][17] ), .A1(\reg_mem[26][17] ), .S(net87544), 
        .Z(n2991) );
  CMXI2X1 U4409 ( .A0(\reg_mem[22][17] ), .A1(\reg_mem[30][17] ), .S(net87520), 
        .Z(n2993) );
  CMXI2X1 U4410 ( .A0(n2994), .A1(n2993), .S(n2190), .Z(n2995) );
  CMXI2X1 U4411 ( .A0(\reg_mem[17][17] ), .A1(\reg_mem[25][17] ), .S(net87545), 
        .Z(n2998) );
  CMXI2X1 U4412 ( .A0(\reg_mem[19][17] ), .A1(\reg_mem[27][17] ), .S(net87525), 
        .Z(n2997) );
  CMXI2X1 U4413 ( .A0(n2998), .A1(n2997), .S(n2181), .Z(n3002) );
  CMXI2X1 U4414 ( .A0(\reg_mem[21][17] ), .A1(\reg_mem[29][17] ), .S(net87524), 
        .Z(n3000) );
  CMXI2X1 U4415 ( .A0(\reg_mem[23][17] ), .A1(\reg_mem[31][17] ), .S(net87522), 
        .Z(n2999) );
  CMXI2X1 U4416 ( .A0(n3002), .A1(n3001), .S(net87248), .Z(n3003) );
  CANR2X1 U4417 ( .A(N185), .B(n3704), .C(N153), .D(n3701), .Z(n3007) );
  CMXI2X1 U4418 ( .A0(\reg_mem[2][16] ), .A1(\reg_mem[10][16] ), .S(net87522), 
        .Z(n3008) );
  CMXI2X1 U4419 ( .A0(n3009), .A1(n3008), .S(n2197), .Z(n3013) );
  CMXI2X1 U4420 ( .A0(\reg_mem[4][16] ), .A1(\reg_mem[12][16] ), .S(net87541), 
        .Z(n3011) );
  CMXI2X1 U4421 ( .A0(\reg_mem[6][16] ), .A1(\reg_mem[14][16] ), .S(net87525), 
        .Z(n3010) );
  CMXI2X1 U4422 ( .A0(n3013), .A1(n3012), .S(n1480), .Z(n3021) );
  CMXI2X1 U4423 ( .A0(\reg_mem[1][16] ), .A1(\reg_mem[9][16] ), .S(net87523), 
        .Z(n3015) );
  CMXI2X1 U4424 ( .A0(\reg_mem[3][16] ), .A1(\reg_mem[11][16] ), .S(net87531), 
        .Z(n3014) );
  CMXI2X1 U4425 ( .A0(n3015), .A1(n3014), .S(n2177), .Z(n3019) );
  CMXI2X1 U4426 ( .A0(\reg_mem[7][16] ), .A1(\reg_mem[15][16] ), .S(net87544), 
        .Z(n3016) );
  CMXI2X1 U4427 ( .A0(n3017), .A1(n3016), .S(n2200), .Z(n3018) );
  CMXI2X1 U4428 ( .A0(n3019), .A1(n3018), .S(net87281), .Z(n3020) );
  CMXI2X1 U4429 ( .A0(n3021), .A1(n3020), .S(net87404), .Z(n3037) );
  CMXI2X1 U4430 ( .A0(\reg_mem[16][16] ), .A1(\reg_mem[24][16] ), .S(net87540), 
        .Z(n3023) );
  CMXI2X1 U4431 ( .A0(\reg_mem[18][16] ), .A1(\reg_mem[26][16] ), .S(net87526), 
        .Z(n3022) );
  CMXI2X1 U4432 ( .A0(\reg_mem[20][16] ), .A1(\reg_mem[28][16] ), .S(net87521), 
        .Z(n3025) );
  CMXI2X1 U4433 ( .A0(\reg_mem[22][16] ), .A1(\reg_mem[30][16] ), .S(net87523), 
        .Z(n3024) );
  CMXI2X1 U4434 ( .A0(n3025), .A1(n3024), .S(n2165), .Z(n3026) );
  CMXI2X1 U4435 ( .A0(n3027), .A1(n3026), .S(net87248), .Z(n3035) );
  CMXI2X1 U4436 ( .A0(\reg_mem[17][16] ), .A1(\reg_mem[25][16] ), .S(net87526), 
        .Z(n3029) );
  CMXI2X1 U4437 ( .A0(\reg_mem[19][16] ), .A1(\reg_mem[27][16] ), .S(net87540), 
        .Z(n3028) );
  CMXI2X1 U4438 ( .A0(\reg_mem[21][16] ), .A1(\reg_mem[29][16] ), .S(net87519), 
        .Z(n3031) );
  CMXI2X1 U4439 ( .A0(n3031), .A1(n3030), .S(n2196), .Z(n3032) );
  CMXI2X1 U4440 ( .A0(n3033), .A1(n3032), .S(net87252), .Z(n3034) );
  CMXI2X1 U4441 ( .A0(n3035), .A1(n3034), .S(net87389), .Z(n3036) );
  CMXI2X1 U4442 ( .A0(n3037), .A1(n3036), .S(n2094), .Z(n3039) );
  CMXI2X1 U4443 ( .A0(n3039), .A1(n3038), .S(n1533), .Z(N285) );
  CIVX2 U4444 ( .A(N111), .Z(n3043) );
  CND2IX1 U4445 ( .B(n3181), .A(N152), .Z(n3042) );
  CIVX2 U4446 ( .A(N79), .Z(n3040) );
  COND3X1 U4447 ( .A(n2115), .B(n3043), .C(n3042), .D(n3041), .Z(n3081) );
  CIVX2 U4448 ( .A(\reg_mem[5][15] ), .Z(n4377) );
  CIVX2 U4449 ( .A(\reg_mem[21][15] ), .Z(n4407) );
  CIVX2 U4450 ( .A(\reg_mem[7][15] ), .Z(n4379) );
  CIVX2 U4451 ( .A(\reg_mem[23][15] ), .Z(n4409) );
  CND2IX1 U4452 ( .B(n3649), .A(n3046), .Z(n3055) );
  CIVX2 U4453 ( .A(\reg_mem[9][15] ), .Z(n4385) );
  CIVX2 U4454 ( .A(\reg_mem[25][15] ), .Z(n4415) );
  CMXI2X1 U4455 ( .A0(n4385), .A1(n4415), .S(n2083), .Z(n3048) );
  CIVX2 U4456 ( .A(\reg_mem[11][15] ), .Z(n4387) );
  CIVX2 U4457 ( .A(\reg_mem[27][15] ), .Z(n4417) );
  CMXI2X1 U4458 ( .A0(n4387), .A1(n4417), .S(n2091), .Z(n3047) );
  CMXI2X1 U4459 ( .A0(n3048), .A1(n3047), .S(n2192), .Z(n3049) );
  CIVX2 U4460 ( .A(\reg_mem[13][15] ), .Z(n4391) );
  CMXI2X1 U4461 ( .A0(n4391), .A1(n4421), .S(n2097), .Z(n3051) );
  CIVX2 U4462 ( .A(\reg_mem[15][15] ), .Z(n4393) );
  CIVX2 U4463 ( .A(\reg_mem[31][15] ), .Z(n4423) );
  CMXI2X1 U4464 ( .A0(n4393), .A1(n4423), .S(n2102), .Z(n3050) );
  CMXI2X1 U4465 ( .A0(n3051), .A1(n3050), .S(n2178), .Z(n3052) );
  CIVX2 U4466 ( .A(\reg_mem[8][15] ), .Z(n4386) );
  CIVX2 U4467 ( .A(\reg_mem[24][15] ), .Z(n4416) );
  CMXI2X1 U4468 ( .A0(n4386), .A1(n4416), .S(n1975), .Z(n3057) );
  CIVX2 U4469 ( .A(\reg_mem[10][15] ), .Z(n4388) );
  CIVX2 U4470 ( .A(\reg_mem[26][15] ), .Z(n4418) );
  CMXI2X1 U4471 ( .A0(n4388), .A1(n4418), .S(n2099), .Z(n3056) );
  CMXI2X1 U4472 ( .A0(n3057), .A1(n3056), .S(n2181), .Z(n3058) );
  CIVX2 U4473 ( .A(\reg_mem[12][15] ), .Z(n4392) );
  CIVX2 U4474 ( .A(\reg_mem[28][15] ), .Z(n4422) );
  CMXI2X1 U4475 ( .A0(n4392), .A1(n4422), .S(n2085), .Z(n3060) );
  CIVX2 U4476 ( .A(\reg_mem[14][15] ), .Z(n4394) );
  CIVX2 U4477 ( .A(\reg_mem[30][15] ), .Z(n4424) );
  CMXI2X1 U4478 ( .A0(n3060), .A1(n3059), .S(n2177), .Z(n3061) );
  CND2IX1 U4479 ( .B(n3667), .A(n3061), .Z(n3066) );
  CIVX2 U4480 ( .A(\reg_mem[1][15] ), .Z(n4371) );
  CIVX2 U4481 ( .A(\reg_mem[17][15] ), .Z(n4401) );
  CMXI2X1 U4482 ( .A0(n4371), .A1(n4401), .S(n2095), .Z(n3063) );
  CIVX2 U4483 ( .A(\reg_mem[3][15] ), .Z(n4373) );
  CIVX2 U4484 ( .A(\reg_mem[19][15] ), .Z(n4403) );
  CMXI2X1 U4485 ( .A0(n4373), .A1(n4403), .S(n2094), .Z(n3062) );
  CMXI2X1 U4486 ( .A0(n3063), .A1(n3062), .S(n2177), .Z(n3064) );
  CND2IX1 U4487 ( .B(n3671), .A(n3064), .Z(n3065) );
  CMXI2X1 U4488 ( .A0(\reg_mem[0][15] ), .A1(\reg_mem[16][15] ), .S(n2101), 
        .Z(n3069) );
  CMXI2X1 U4489 ( .A0(\reg_mem[2][15] ), .A1(\reg_mem[18][15] ), .S(n2084), 
        .Z(n3068) );
  CMXI2X1 U4490 ( .A0(n3069), .A1(n3068), .S(n2200), .Z(n3073) );
  CMXI2X1 U4491 ( .A0(\reg_mem[4][15] ), .A1(\reg_mem[20][15] ), .S(n2089), 
        .Z(n3071) );
  CMXI2X1 U4492 ( .A0(n3071), .A1(n3070), .S(n2179), .Z(n3072) );
  CIVX2 U4493 ( .A(N110), .Z(n3084) );
  CND2IX1 U4494 ( .B(n3181), .A(N151), .Z(n3082) );
  CMXI2X1 U4495 ( .A0(\reg_mem[0][14] ), .A1(\reg_mem[8][14] ), .S(net87522), 
        .Z(n3088) );
  CMXI2X1 U4496 ( .A0(\reg_mem[2][14] ), .A1(\reg_mem[10][14] ), .S(net87523), 
        .Z(n3087) );
  CMXI2X1 U4497 ( .A0(\reg_mem[4][14] ), .A1(\reg_mem[12][14] ), .S(net87524), 
        .Z(n3090) );
  CMXI2X1 U4498 ( .A0(\reg_mem[6][14] ), .A1(\reg_mem[14][14] ), .S(net87533), 
        .Z(n3089) );
  CMXI2X1 U4499 ( .A0(n3092), .A1(n3091), .S(net87262), .Z(n3100) );
  CMXI2X1 U4500 ( .A0(\reg_mem[1][14] ), .A1(\reg_mem[9][14] ), .S(net87525), 
        .Z(n3094) );
  CMXI2X1 U4501 ( .A0(\reg_mem[3][14] ), .A1(\reg_mem[11][14] ), .S(net87526), 
        .Z(n3093) );
  CMXI2X1 U4502 ( .A0(\reg_mem[7][14] ), .A1(\reg_mem[15][14] ), .S(net87529), 
        .Z(n3095) );
  CMXI2X1 U4503 ( .A0(n3098), .A1(n3097), .S(net87279), .Z(n3099) );
  CMXI2X1 U4504 ( .A0(\reg_mem[16][14] ), .A1(\reg_mem[24][14] ), .S(net87532), 
        .Z(n3102) );
  CMXI2X1 U4505 ( .A0(\reg_mem[18][14] ), .A1(\reg_mem[26][14] ), .S(net87532), 
        .Z(n3101) );
  CMXI2X1 U4506 ( .A0(\reg_mem[20][14] ), .A1(\reg_mem[28][14] ), .S(net87531), 
        .Z(n3104) );
  CMXI2X1 U4507 ( .A0(\reg_mem[22][14] ), .A1(\reg_mem[30][14] ), .S(net87519), 
        .Z(n3103) );
  CMXI2X1 U4508 ( .A0(\reg_mem[17][14] ), .A1(\reg_mem[25][14] ), .S(net87538), 
        .Z(n3108) );
  CMXI2X1 U4509 ( .A0(\reg_mem[19][14] ), .A1(\reg_mem[27][14] ), .S(net87522), 
        .Z(n3107) );
  CMXI2X1 U4510 ( .A0(\reg_mem[23][14] ), .A1(\reg_mem[31][14] ), .S(net87525), 
        .Z(n3109) );
  CIVX2 U4511 ( .A(N109), .Z(n3117) );
  CIVX2 U4512 ( .A(N77), .Z(n3115) );
  CANR2X1 U4513 ( .A(N182), .B(n3704), .C(N150), .D(n3701), .Z(n3118) );
  CMXI2X1 U4514 ( .A0(net79481), .A1(net79482), .S(n2196), .Z(n3123) );
  CMXI2X1 U4515 ( .A0(\reg_mem[4][13] ), .A1(\reg_mem[12][13] ), .S(net87529), 
        .Z(n3121) );
  CMXI2X1 U4516 ( .A0(n3121), .A1(n3120), .S(n2183), .Z(n3122) );
  CMXI2X1 U4517 ( .A0(n3123), .A1(n3122), .S(net87261), .Z(n3129) );
  CMXI2X1 U4518 ( .A0(net79475), .A1(net79476), .S(n2166), .Z(n3127) );
  CMXI2X1 U4519 ( .A0(\reg_mem[5][13] ), .A1(\reg_mem[13][13] ), .S(net87530), 
        .Z(n3125) );
  CMXI2X1 U4520 ( .A0(\reg_mem[7][13] ), .A1(\reg_mem[15][13] ), .S(net87524), 
        .Z(n3124) );
  CMXI2X1 U4521 ( .A0(n3127), .A1(n3126), .S(net87275), .Z(n3128) );
  CMXI2X1 U4522 ( .A0(n3129), .A1(n3128), .S(net87401), .Z(n3144) );
  CMXI2X1 U4523 ( .A0(\reg_mem[16][13] ), .A1(\reg_mem[20][13] ), .S(net87251), 
        .Z(n3131) );
  CMXI2X1 U4524 ( .A0(\reg_mem[18][13] ), .A1(\reg_mem[22][13] ), .S(net87277), 
        .Z(n3130) );
  CMXI2X1 U4525 ( .A0(n3131), .A1(n3130), .S(n2192), .Z(n3135) );
  CMXI2X1 U4526 ( .A0(\reg_mem[17][13] ), .A1(\reg_mem[21][13] ), .S(net87253), 
        .Z(n3133) );
  CMXI2X1 U4527 ( .A0(\reg_mem[19][13] ), .A1(\reg_mem[23][13] ), .S(net87255), 
        .Z(n3132) );
  CMXI2X1 U4528 ( .A0(n3133), .A1(n3132), .S(n2165), .Z(n3134) );
  CMXI2X1 U4529 ( .A0(\reg_mem[24][13] ), .A1(\reg_mem[28][13] ), .S(net87277), 
        .Z(n3137) );
  CMXI2X1 U4530 ( .A0(\reg_mem[26][13] ), .A1(\reg_mem[30][13] ), .S(net87256), 
        .Z(n3136) );
  CMXI2X1 U4531 ( .A0(n3137), .A1(n3136), .S(n1469), .Z(n3141) );
  CMXI2X1 U4532 ( .A0(\reg_mem[25][13] ), .A1(\reg_mem[29][13] ), .S(net87260), 
        .Z(n3139) );
  CMXI2X1 U4533 ( .A0(\reg_mem[27][13] ), .A1(\reg_mem[31][13] ), .S(net87266), 
        .Z(n3138) );
  CMXI2X1 U4534 ( .A0(n3139), .A1(n3138), .S(n2165), .Z(n3140) );
  CMXI2X1 U4535 ( .A0(n3141), .A1(n3140), .S(net87403), .Z(n3142) );
  CANR2X1 U4536 ( .A(N181), .B(n3704), .C(N149), .D(n3701), .Z(n3148) );
  CMXI2X1 U4537 ( .A0(\reg_mem[0][12] ), .A1(\reg_mem[4][12] ), .S(net87255), 
        .Z(n3150) );
  CMXI2X1 U4538 ( .A0(\reg_mem[2][12] ), .A1(\reg_mem[6][12] ), .S(net87276), 
        .Z(n3149) );
  CMXI2X1 U4539 ( .A0(n3150), .A1(n3149), .S(n2195), .Z(n3154) );
  CMXI2X1 U4540 ( .A0(\reg_mem[1][12] ), .A1(\reg_mem[5][12] ), .S(net87256), 
        .Z(n3152) );
  CMXI2X1 U4541 ( .A0(\reg_mem[3][12] ), .A1(\reg_mem[7][12] ), .S(net87247), 
        .Z(n3151) );
  CMXI2X1 U4542 ( .A0(n3152), .A1(n3151), .S(n2182), .Z(n3153) );
  CMXI2X1 U4543 ( .A0(n3154), .A1(n3153), .S(net87388), .Z(n3162) );
  CMXI2X1 U4544 ( .A0(\reg_mem[8][12] ), .A1(\reg_mem[12][12] ), .S(net87281), 
        .Z(n3156) );
  CMXI2X1 U4545 ( .A0(\reg_mem[10][12] ), .A1(\reg_mem[14][12] ), .S(net87253), 
        .Z(n3155) );
  CMXI2X1 U4546 ( .A0(n3156), .A1(n3155), .S(n2162), .Z(n3160) );
  CMXI2X1 U4547 ( .A0(\reg_mem[9][12] ), .A1(\reg_mem[13][12] ), .S(net87261), 
        .Z(n3158) );
  CMXI2X1 U4548 ( .A0(\reg_mem[11][12] ), .A1(\reg_mem[15][12] ), .S(net87273), 
        .Z(n3157) );
  CMXI2X1 U4549 ( .A0(n3160), .A1(n3159), .S(net87389), .Z(n3161) );
  CMXI2X1 U4550 ( .A0(\reg_mem[16][12] ), .A1(\reg_mem[20][12] ), .S(net87242), 
        .Z(n3164) );
  CMXI2X1 U4551 ( .A0(\reg_mem[18][12] ), .A1(\reg_mem[22][12] ), .S(net87258), 
        .Z(n3163) );
  CMXI2X1 U4552 ( .A0(n3164), .A1(n3163), .S(n2191), .Z(n3168) );
  CMXI2X1 U4553 ( .A0(\reg_mem[17][12] ), .A1(\reg_mem[21][12] ), .S(net87268), 
        .Z(n3166) );
  CMXI2X1 U4554 ( .A0(\reg_mem[19][12] ), .A1(\reg_mem[23][12] ), .S(net87271), 
        .Z(n3165) );
  CMXI2X1 U4555 ( .A0(n3168), .A1(n3167), .S(net87392), .Z(n3176) );
  CMXI2X1 U4556 ( .A0(\reg_mem[26][12] ), .A1(\reg_mem[30][12] ), .S(net87263), 
        .Z(n3169) );
  CMXI2X1 U4557 ( .A0(\reg_mem[25][12] ), .A1(\reg_mem[29][12] ), .S(net87269), 
        .Z(n3172) );
  CMXI2X1 U4558 ( .A0(\reg_mem[27][12] ), .A1(\reg_mem[31][12] ), .S(net87265), 
        .Z(n3171) );
  CMXI2X1 U4559 ( .A0(n3172), .A1(n3171), .S(n2195), .Z(n3173) );
  CMXI2X1 U4560 ( .A0(n3174), .A1(n3173), .S(net87863), .Z(n3175) );
  CMXI2X1 U4561 ( .A0(n3176), .A1(n3175), .S(n1532), .Z(n3177) );
  CIVX2 U4562 ( .A(alu_op_c[12]), .Z(n3179) );
  CIVX2 U4563 ( .A(N107), .Z(n3184) );
  CND2IX1 U4564 ( .B(n3181), .A(N148), .Z(n3182) );
  CND2IX1 U4565 ( .B(n3186), .A(n3185), .Z(alu_op_c[11]) );
  CMXI2X1 U4566 ( .A0(net79408), .A1(net79409), .S(n2194), .Z(n3188) );
  CMXI2X1 U4567 ( .A0(net79406), .A1(net79407), .S(n2181), .Z(n3187) );
  CMXI2X1 U4568 ( .A0(n3188), .A1(n3187), .S(net87410), .Z(n3196) );
  CMXI2X1 U4569 ( .A0(\reg_mem[8][11] ), .A1(\reg_mem[12][11] ), .S(net87281), 
        .Z(n3190) );
  CMXI2X1 U4570 ( .A0(\reg_mem[10][11] ), .A1(\reg_mem[14][11] ), .S(net87263), 
        .Z(n3189) );
  CMXI2X1 U4571 ( .A0(\reg_mem[9][11] ), .A1(\reg_mem[13][11] ), .S(net87272), 
        .Z(n3192) );
  CMXI2X1 U4572 ( .A0(\reg_mem[11][11] ), .A1(\reg_mem[15][11] ), .S(net87277), 
        .Z(n3191) );
  CMXI2X1 U4573 ( .A0(n3192), .A1(n3191), .S(n2162), .Z(n3193) );
  CMXI2X1 U4574 ( .A0(\reg_mem[16][11] ), .A1(\reg_mem[17][11] ), .S(net87406), 
        .Z(n3198) );
  CMXI2X1 U4575 ( .A0(n3198), .A1(n3197), .S(n2190), .Z(n3202) );
  CMXI2X1 U4576 ( .A0(\reg_mem[20][11] ), .A1(\reg_mem[21][11] ), .S(net87393), 
        .Z(n3200) );
  CMXI2X1 U4577 ( .A0(\reg_mem[22][11] ), .A1(\reg_mem[23][11] ), .S(net87393), 
        .Z(n3199) );
  CMXI2X1 U4578 ( .A0(n3200), .A1(n3199), .S(n2186), .Z(n3201) );
  CMXI2X1 U4579 ( .A0(n3202), .A1(n3201), .S(net87279), .Z(n3210) );
  CMXI2X1 U4580 ( .A0(\reg_mem[24][11] ), .A1(\reg_mem[25][11] ), .S(n2069), 
        .Z(n3204) );
  CMXI2X1 U4581 ( .A0(\reg_mem[26][11] ), .A1(\reg_mem[27][11] ), .S(net87403), 
        .Z(n3203) );
  CMXI2X1 U4582 ( .A0(n3204), .A1(n3203), .S(n2179), .Z(n3208) );
  CMXI2X1 U4583 ( .A0(\reg_mem[28][11] ), .A1(\reg_mem[29][11] ), .S(net87397), 
        .Z(n3206) );
  CMXI2X1 U4584 ( .A0(\reg_mem[30][11] ), .A1(\reg_mem[31][11] ), .S(net87411), 
        .Z(n3205) );
  CMXI2X1 U4585 ( .A0(n3206), .A1(n3205), .S(n2194), .Z(n3207) );
  CMXI2X1 U4586 ( .A0(n3208), .A1(n3207), .S(net87248), .Z(n3209) );
  CMXI2X1 U4587 ( .A0(n3210), .A1(n3209), .S(net87533), .Z(n3211) );
  CANR2X1 U4588 ( .A(N179), .B(n3704), .C(N147), .D(n3701), .Z(n3217) );
  CMXI2X1 U4589 ( .A0(\reg_mem[0][10] ), .A1(\reg_mem[1][10] ), .S(net87393), 
        .Z(n3219) );
  CMXI2X1 U4590 ( .A0(\reg_mem[2][10] ), .A1(\reg_mem[3][10] ), .S(net87389), 
        .Z(n3218) );
  CMXI2X1 U4591 ( .A0(n3219), .A1(n3218), .S(n2197), .Z(n3223) );
  CMXI2X1 U4592 ( .A0(\reg_mem[4][10] ), .A1(\reg_mem[5][10] ), .S(net87412), 
        .Z(n3221) );
  CMXI2X1 U4593 ( .A0(\reg_mem[6][10] ), .A1(\reg_mem[7][10] ), .S(net87399), 
        .Z(n3220) );
  CMXI2X1 U4594 ( .A0(n3221), .A1(n3220), .S(n2193), .Z(n3222) );
  CMXI2X1 U4595 ( .A0(n3223), .A1(n3222), .S(n1391), .Z(n3231) );
  CMXI2X1 U4596 ( .A0(\reg_mem[8][10] ), .A1(\reg_mem[9][10] ), .S(n1456), .Z(
        n3225) );
  CMXI2X1 U4597 ( .A0(\reg_mem[10][10] ), .A1(\reg_mem[11][10] ), .S(net87412), 
        .Z(n3224) );
  CMXI2X1 U4598 ( .A0(n3225), .A1(n3224), .S(n2179), .Z(n3229) );
  CMXI2X1 U4599 ( .A0(\reg_mem[12][10] ), .A1(\reg_mem[13][10] ), .S(net87402), 
        .Z(n3227) );
  CMXI2X1 U4600 ( .A0(\reg_mem[14][10] ), .A1(\reg_mem[15][10] ), .S(net87385), 
        .Z(n3226) );
  CMXI2X1 U4601 ( .A0(n3227), .A1(n3226), .S(n2179), .Z(n3228) );
  CMXI2X1 U4602 ( .A0(n3229), .A1(n3228), .S(net87267), .Z(n3230) );
  CMXI2X1 U4603 ( .A0(n3231), .A1(n3230), .S(net87856), .Z(n3247) );
  CMXI2X1 U4604 ( .A0(\reg_mem[16][10] ), .A1(\reg_mem[17][10] ), .S(net87402), 
        .Z(n3233) );
  CMXI2X1 U4605 ( .A0(\reg_mem[18][10] ), .A1(\reg_mem[19][10] ), .S(net87408), 
        .Z(n3232) );
  CMXI2X1 U4606 ( .A0(n3233), .A1(n3232), .S(n2185), .Z(n3237) );
  CMXI2X1 U4607 ( .A0(\reg_mem[20][10] ), .A1(\reg_mem[21][10] ), .S(net87387), 
        .Z(n3235) );
  CMXI2X1 U4608 ( .A0(\reg_mem[22][10] ), .A1(\reg_mem[23][10] ), .S(net87389), 
        .Z(n3234) );
  CMXI2X1 U4609 ( .A0(n3235), .A1(n3234), .S(n2186), .Z(n3236) );
  CMXI2X1 U4610 ( .A0(n3237), .A1(n3236), .S(net87280), .Z(n3245) );
  CMXI2X1 U4611 ( .A0(\reg_mem[24][10] ), .A1(\reg_mem[25][10] ), .S(net87387), 
        .Z(n3239) );
  CMXI2X1 U4612 ( .A0(\reg_mem[26][10] ), .A1(\reg_mem[27][10] ), .S(net87395), 
        .Z(n3238) );
  CMXI2X1 U4613 ( .A0(\reg_mem[28][10] ), .A1(\reg_mem[29][10] ), .S(net87404), 
        .Z(n3241) );
  CMXI2X1 U4614 ( .A0(\reg_mem[30][10] ), .A1(\reg_mem[31][10] ), .S(net87404), 
        .Z(n3240) );
  CMXI2X1 U4615 ( .A0(n3241), .A1(n3240), .S(n2193), .Z(n3242) );
  CMXI2X1 U4616 ( .A0(n3243), .A1(n3242), .S(n1385), .Z(n3244) );
  CANR2X1 U4617 ( .A(N178), .B(n3704), .C(N146), .D(n3701), .Z(n3252) );
  CMXI2X1 U4618 ( .A0(\reg_mem[0][9] ), .A1(\reg_mem[1][9] ), .S(net87403), 
        .Z(n3254) );
  CMXI2X1 U4619 ( .A0(\reg_mem[2][9] ), .A1(\reg_mem[3][9] ), .S(net87411), 
        .Z(n3253) );
  CMXI2X1 U4620 ( .A0(n3254), .A1(n3253), .S(n2196), .Z(n3258) );
  CMXI2X1 U4621 ( .A0(\reg_mem[4][9] ), .A1(\reg_mem[5][9] ), .S(net87406), 
        .Z(n3256) );
  CMXI2X1 U4622 ( .A0(\reg_mem[6][9] ), .A1(\reg_mem[7][9] ), .S(net87394), 
        .Z(n3255) );
  CMXI2X1 U4623 ( .A0(n3256), .A1(n3255), .S(n2192), .Z(n3257) );
  CMXI2X1 U4624 ( .A0(n3258), .A1(n3257), .S(net87247), .Z(n3266) );
  CMXI2X1 U4625 ( .A0(\reg_mem[10][9] ), .A1(\reg_mem[11][9] ), .S(net87398), 
        .Z(n3259) );
  CMXI2X1 U4626 ( .A0(n3260), .A1(n3259), .S(n2178), .Z(n3264) );
  CMXI2X1 U4627 ( .A0(\reg_mem[12][9] ), .A1(\reg_mem[13][9] ), .S(net87388), 
        .Z(n3262) );
  CMXI2X1 U4628 ( .A0(\reg_mem[14][9] ), .A1(\reg_mem[15][9] ), .S(net87397), 
        .Z(n3261) );
  CMXI2X1 U4629 ( .A0(n3262), .A1(n3261), .S(n2178), .Z(n3263) );
  CMXI2X1 U4630 ( .A0(n3264), .A1(n3263), .S(net87260), .Z(n3265) );
  CMXI2X1 U4631 ( .A0(n3266), .A1(n3265), .S(n1532), .Z(n3282) );
  CMXI2X1 U4632 ( .A0(\reg_mem[16][9] ), .A1(\reg_mem[17][9] ), .S(net87385), 
        .Z(n3268) );
  CMXI2X1 U4633 ( .A0(\reg_mem[18][9] ), .A1(\reg_mem[19][9] ), .S(net87401), 
        .Z(n3267) );
  CMXI2X1 U4634 ( .A0(n3268), .A1(n3267), .S(n2184), .Z(n3272) );
  CMXI2X1 U4635 ( .A0(\reg_mem[20][9] ), .A1(\reg_mem[21][9] ), .S(net87386), 
        .Z(n3270) );
  CMXI2X1 U4636 ( .A0(\reg_mem[22][9] ), .A1(\reg_mem[23][9] ), .S(net87392), 
        .Z(n3269) );
  CMXI2X1 U4637 ( .A0(n3270), .A1(n3269), .S(n2185), .Z(n3271) );
  CMXI2X1 U4638 ( .A0(n3272), .A1(n3271), .S(n1480), .Z(n3280) );
  CMXI2X1 U4639 ( .A0(\reg_mem[24][9] ), .A1(\reg_mem[25][9] ), .S(net87402), 
        .Z(n3274) );
  CMXI2X1 U4640 ( .A0(\reg_mem[26][9] ), .A1(\reg_mem[27][9] ), .S(net87404), 
        .Z(n3273) );
  CMXI2X1 U4641 ( .A0(\reg_mem[28][9] ), .A1(\reg_mem[29][9] ), .S(net87403), 
        .Z(n3276) );
  CMXI2X1 U4642 ( .A0(\reg_mem[30][9] ), .A1(\reg_mem[31][9] ), .S(net87408), 
        .Z(n3275) );
  CMXI2X1 U4643 ( .A0(n3280), .A1(n3279), .S(net87856), .Z(n3281) );
  CIVX2 U4644 ( .A(alu_op_c[9]), .Z(n3283) );
  CANR2X1 U4645 ( .A(N144), .B(n3701), .C(n3476), .D(n3285), .Z(n3290) );
  CMXI2X1 U4646 ( .A0(\reg_mem[0][7] ), .A1(\reg_mem[1][7] ), .S(net87412), 
        .Z(n3292) );
  CMXI2X1 U4647 ( .A0(\reg_mem[2][7] ), .A1(\reg_mem[3][7] ), .S(net87412), 
        .Z(n3291) );
  CMXI2X1 U4648 ( .A0(n3292), .A1(n3291), .S(n2199), .Z(n3296) );
  CMXI2X1 U4649 ( .A0(\reg_mem[6][7] ), .A1(\reg_mem[7][7] ), .S(net87398), 
        .Z(n3293) );
  CMXI2X1 U4650 ( .A0(n3294), .A1(n3293), .S(n2191), .Z(n3295) );
  CMXI2X1 U4651 ( .A0(n3296), .A1(n3295), .S(net87253), .Z(n3304) );
  CMXI2X1 U4652 ( .A0(\reg_mem[8][7] ), .A1(\reg_mem[9][7] ), .S(net87410), 
        .Z(n3298) );
  CMXI2X1 U4653 ( .A0(\reg_mem[10][7] ), .A1(\reg_mem[11][7] ), .S(net87386), 
        .Z(n3297) );
  CMXI2X1 U4654 ( .A0(n3298), .A1(n3297), .S(n2180), .Z(n3302) );
  CMXI2X1 U4655 ( .A0(\reg_mem[12][7] ), .A1(\reg_mem[13][7] ), .S(net87397), 
        .Z(n3300) );
  CMXI2X1 U4656 ( .A0(\reg_mem[14][7] ), .A1(\reg_mem[15][7] ), .S(n2070), .Z(
        n3299) );
  CMXI2X1 U4657 ( .A0(n3300), .A1(n3299), .S(n2165), .Z(n3301) );
  CMXI2X1 U4658 ( .A0(n3302), .A1(n3301), .S(net87262), .Z(n3303) );
  CMXI2X1 U4659 ( .A0(n3304), .A1(n3303), .S(n1460), .Z(n3320) );
  CMXI2X1 U4660 ( .A0(\reg_mem[16][7] ), .A1(\reg_mem[17][7] ), .S(n1456), .Z(
        n3306) );
  CMXI2X1 U4661 ( .A0(\reg_mem[18][7] ), .A1(\reg_mem[19][7] ), .S(net87388), 
        .Z(n3305) );
  CMXI2X1 U4662 ( .A0(n3306), .A1(n3305), .S(n2165), .Z(n3310) );
  CMXI2X1 U4663 ( .A0(\reg_mem[20][7] ), .A1(\reg_mem[21][7] ), .S(net87410), 
        .Z(n3308) );
  CMXI2X1 U4664 ( .A0(\reg_mem[22][7] ), .A1(\reg_mem[23][7] ), .S(net87385), 
        .Z(n3307) );
  CMXI2X1 U4665 ( .A0(n3308), .A1(n3307), .S(n2189), .Z(n3309) );
  CMXI2X1 U4666 ( .A0(n3310), .A1(n3309), .S(net87266), .Z(n3318) );
  CMXI2X1 U4667 ( .A0(\reg_mem[24][7] ), .A1(\reg_mem[25][7] ), .S(net87385), 
        .Z(n3312) );
  CMXI2X1 U4668 ( .A0(\reg_mem[26][7] ), .A1(\reg_mem[27][7] ), .S(n1456), .Z(
        n3311) );
  CMXI2X1 U4669 ( .A0(n3312), .A1(n3311), .S(n2200), .Z(n3316) );
  CMXI2X1 U4670 ( .A0(\reg_mem[28][7] ), .A1(\reg_mem[29][7] ), .S(net87385), 
        .Z(n3314) );
  CMXI2X1 U4671 ( .A0(\reg_mem[30][7] ), .A1(\reg_mem[31][7] ), .S(net87391), 
        .Z(n3313) );
  CMXI2X1 U4672 ( .A0(n3314), .A1(n3313), .S(n2195), .Z(n3315) );
  CMXI2X1 U4673 ( .A0(n3316), .A1(n3315), .S(n1480), .Z(n3317) );
  CMXI2X1 U4674 ( .A0(n3318), .A1(n3317), .S(net87540), .Z(n3319) );
  CMXI2X1 U4675 ( .A0(n3320), .A1(n3319), .S(n2099), .Z(n3322) );
  CIVX2 U4676 ( .A(alu_op_c[7]), .Z(n3321) );
  CENX1 U4677 ( .A(prog_count_ex[6]), .B(n3382), .Z(n3323) );
  CANR2X1 U4678 ( .A(N143), .B(n3701), .C(n3476), .D(n3323), .Z(n3324) );
  CIVX2 U4679 ( .A(n3324), .Z(n3325) );
  CIVX2 U4680 ( .A(opcode_ext_ex[1]), .Z(n3342) );
  CND2IX1 U4681 ( .B(opcode_ex[2]), .A(opcode_ex[5]), .Z(n3331) );
  CIVX2 U4682 ( .A(n3331), .Z(n5238) );
  CND2IX1 U4683 ( .B(opcode_ext_ex[10]), .A(n3335), .Z(n3338) );
  CND2IX1 U4684 ( .B(opcode_ext_ex[7]), .A(n3336), .Z(n3337) );
  CIVX2 U4685 ( .A(n3437), .Z(n3750) );
  CIVX2 U4686 ( .A(n3751), .Z(n3739) );
  CMXI2X1 U4687 ( .A0(\reg_mem[0][6] ), .A1(\reg_mem[1][6] ), .S(n2070), .Z(
        n3350) );
  CMXI2X1 U4688 ( .A0(\reg_mem[2][6] ), .A1(\reg_mem[3][6] ), .S(net87399), 
        .Z(n3349) );
  CMXI2X1 U4689 ( .A0(n3350), .A1(n3349), .S(n2200), .Z(n3354) );
  CMXI2X1 U4690 ( .A0(\reg_mem[4][6] ), .A1(\reg_mem[5][6] ), .S(net87395), 
        .Z(n3352) );
  CMXI2X1 U4691 ( .A0(\reg_mem[6][6] ), .A1(\reg_mem[7][6] ), .S(net87392), 
        .Z(n3351) );
  CMXI2X1 U4692 ( .A0(n3352), .A1(n3351), .S(n2194), .Z(n3353) );
  CMXI2X1 U4693 ( .A0(n3354), .A1(n3353), .S(net87248), .Z(n3362) );
  CMXI2X1 U4694 ( .A0(\reg_mem[8][6] ), .A1(\reg_mem[9][6] ), .S(net87385), 
        .Z(n3356) );
  CMXI2X1 U4695 ( .A0(\reg_mem[10][6] ), .A1(\reg_mem[11][6] ), .S(net87396), 
        .Z(n3355) );
  CMXI2X1 U4696 ( .A0(n3356), .A1(n3355), .S(n2180), .Z(n3360) );
  CMXI2X1 U4697 ( .A0(\reg_mem[12][6] ), .A1(\reg_mem[13][6] ), .S(net87387), 
        .Z(n3358) );
  CMXI2X1 U4698 ( .A0(\reg_mem[14][6] ), .A1(\reg_mem[15][6] ), .S(net87397), 
        .Z(n3357) );
  CMXI2X1 U4699 ( .A0(n3358), .A1(n3357), .S(n2180), .Z(n3359) );
  CMXI2X1 U4700 ( .A0(n3360), .A1(n3359), .S(net87253), .Z(n3361) );
  CMXI2X1 U4701 ( .A0(n3362), .A1(n3361), .S(net87544), .Z(n3378) );
  CMXI2X1 U4702 ( .A0(\reg_mem[16][6] ), .A1(\reg_mem[17][6] ), .S(net87386), 
        .Z(n3364) );
  CMXI2X1 U4703 ( .A0(\reg_mem[18][6] ), .A1(\reg_mem[19][6] ), .S(n2069), .Z(
        n3363) );
  CMXI2X1 U4704 ( .A0(n3364), .A1(n3363), .S(n2186), .Z(n3368) );
  CMXI2X1 U4705 ( .A0(\reg_mem[20][6] ), .A1(\reg_mem[21][6] ), .S(net87391), 
        .Z(n3366) );
  CMXI2X1 U4706 ( .A0(\reg_mem[22][6] ), .A1(\reg_mem[23][6] ), .S(net87387), 
        .Z(n3365) );
  CMXI2X1 U4707 ( .A0(n3366), .A1(n3365), .S(n2187), .Z(n3367) );
  CMXI2X1 U4708 ( .A0(n3368), .A1(n3367), .S(net87256), .Z(n3376) );
  CMXI2X1 U4709 ( .A0(\reg_mem[24][6] ), .A1(\reg_mem[25][6] ), .S(net87402), 
        .Z(n3370) );
  CMXI2X1 U4710 ( .A0(\reg_mem[26][6] ), .A1(\reg_mem[27][6] ), .S(net87398), 
        .Z(n3369) );
  CMXI2X1 U4711 ( .A0(n3370), .A1(n3369), .S(n2199), .Z(n3374) );
  CMXI2X1 U4712 ( .A0(\reg_mem[28][6] ), .A1(\reg_mem[29][6] ), .S(net87406), 
        .Z(n3372) );
  CMXI2X1 U4713 ( .A0(\reg_mem[30][6] ), .A1(\reg_mem[31][6] ), .S(net87393), 
        .Z(n3371) );
  CMXI2X1 U4714 ( .A0(n3372), .A1(n3371), .S(n2194), .Z(n3373) );
  CMXI2X1 U4715 ( .A0(n3374), .A1(n3373), .S(net87276), .Z(n3375) );
  CMXI2X1 U4716 ( .A0(n3376), .A1(n3375), .S(net87541), .Z(n3377) );
  CIVX2 U4717 ( .A(N101), .Z(n3391) );
  CIVX2 U4718 ( .A(N69), .Z(n3381) );
  CIVX2 U4719 ( .A(n3384), .Z(n3385) );
  CANR2X1 U4720 ( .A(N142), .B(n3701), .C(n3386), .D(n3385), .Z(n3387) );
  CIVX2 U4721 ( .A(n3387), .Z(n3388) );
  CMXI2X1 U4722 ( .A0(n3393), .A1(n3392), .S(prog_count_o[5]), .Z(n3395) );
  CMXI2X1 U4723 ( .A0(\reg_mem[0][5] ), .A1(\reg_mem[1][5] ), .S(net87399), 
        .Z(n3398) );
  CMXI2X1 U4724 ( .A0(\reg_mem[2][5] ), .A1(\reg_mem[3][5] ), .S(n1456), .Z(
        n3397) );
  CMXI2X1 U4725 ( .A0(n3398), .A1(n3397), .S(n2198), .Z(n3402) );
  CMXI2X1 U4726 ( .A0(\reg_mem[4][5] ), .A1(\reg_mem[5][5] ), .S(net87409), 
        .Z(n3400) );
  CMXI2X1 U4727 ( .A0(\reg_mem[6][5] ), .A1(\reg_mem[7][5] ), .S(net87408), 
        .Z(n3399) );
  CMXI2X1 U4728 ( .A0(n3400), .A1(n3399), .S(n2190), .Z(n3401) );
  CMXI2X1 U4729 ( .A0(\reg_mem[8][5] ), .A1(\reg_mem[9][5] ), .S(net87406), 
        .Z(n3404) );
  CMXI2X1 U4730 ( .A0(\reg_mem[10][5] ), .A1(\reg_mem[11][5] ), .S(net87398), 
        .Z(n3403) );
  CMXI2X1 U4731 ( .A0(\reg_mem[12][5] ), .A1(\reg_mem[13][5] ), .S(net87407), 
        .Z(n3406) );
  CMXI2X1 U4732 ( .A0(\reg_mem[14][5] ), .A1(\reg_mem[15][5] ), .S(net87401), 
        .Z(n3405) );
  CMXI2X1 U4733 ( .A0(n3406), .A1(n3405), .S(n2162), .Z(n3407) );
  CMXI2X1 U4734 ( .A0(\reg_mem[16][5] ), .A1(\reg_mem[17][5] ), .S(net87407), 
        .Z(n3412) );
  CMXI2X1 U4735 ( .A0(\reg_mem[18][5] ), .A1(\reg_mem[19][5] ), .S(net87389), 
        .Z(n3411) );
  CMXI2X1 U4736 ( .A0(n3412), .A1(n3411), .S(n2183), .Z(n3416) );
  CMXI2X1 U4737 ( .A0(\reg_mem[20][5] ), .A1(\reg_mem[21][5] ), .S(net87385), 
        .Z(n3414) );
  CMXI2X1 U4738 ( .A0(\reg_mem[22][5] ), .A1(\reg_mem[23][5] ), .S(net87385), 
        .Z(n3413) );
  CMXI2X1 U4739 ( .A0(n3414), .A1(n3413), .S(n2184), .Z(n3415) );
  CMXI2X1 U4740 ( .A0(n3416), .A1(n3415), .S(net87279), .Z(n3424) );
  CMXI2X1 U4741 ( .A0(\reg_mem[24][5] ), .A1(\reg_mem[25][5] ), .S(net87391), 
        .Z(n3418) );
  CMXI2X1 U4742 ( .A0(\reg_mem[26][5] ), .A1(\reg_mem[27][5] ), .S(net87396), 
        .Z(n3417) );
  CMXI2X1 U4743 ( .A0(\reg_mem[28][5] ), .A1(\reg_mem[29][5] ), .S(net87407), 
        .Z(n3420) );
  CMXI2X1 U4744 ( .A0(\reg_mem[30][5] ), .A1(\reg_mem[31][5] ), .S(net87397), 
        .Z(n3419) );
  CIVX2 U4745 ( .A(alu_op_c[5]), .Z(n3427) );
  CIVX2 U4746 ( .A(N100), .Z(n3436) );
  CIVX2 U4747 ( .A(N68), .Z(n3429) );
  CENX1 U4748 ( .A(prog_count_ex[4]), .B(n3430), .Z(n3431) );
  CANR2X1 U4749 ( .A(N141), .B(n3701), .C(n3476), .D(n3431), .Z(n3432) );
  CIVX2 U4750 ( .A(n3432), .Z(n3433) );
  COND3X1 U4751 ( .A(n2272), .B(n3436), .C(n3435), .D(n3434), .Z(alu_op_c[4])
         );
  CND2IX1 U4752 ( .B(n3437), .A(alu_op_c[4]), .Z(n3443) );
  CND2IX1 U4753 ( .B(n2062), .A(n2146), .Z(n3442) );
  CMXI2X1 U4754 ( .A0(\reg_mem[0][4] ), .A1(\reg_mem[1][4] ), .S(net87400), 
        .Z(n3445) );
  CMXI2X1 U4755 ( .A0(\reg_mem[2][4] ), .A1(\reg_mem[3][4] ), .S(net87389), 
        .Z(n3444) );
  CMXI2X1 U4756 ( .A0(n3445), .A1(n3444), .S(n2197), .Z(n3449) );
  CMXI2X1 U4757 ( .A0(\reg_mem[4][4] ), .A1(\reg_mem[5][4] ), .S(net87410), 
        .Z(n3447) );
  CMXI2X1 U4758 ( .A0(\reg_mem[6][4] ), .A1(\reg_mem[7][4] ), .S(n1456), .Z(
        n3446) );
  CMXI2X1 U4759 ( .A0(n3447), .A1(n3446), .S(n2183), .Z(n3448) );
  CMXI2X1 U4760 ( .A0(n3449), .A1(n3448), .S(net87278), .Z(n3457) );
  CMXI2X1 U4761 ( .A0(\reg_mem[8][4] ), .A1(\reg_mem[9][4] ), .S(net87389), 
        .Z(n3451) );
  CMXI2X1 U4762 ( .A0(\reg_mem[10][4] ), .A1(\reg_mem[11][4] ), .S(net87396), 
        .Z(n3450) );
  CMXI2X1 U4763 ( .A0(n3451), .A1(n3450), .S(n2162), .Z(n3455) );
  CMXI2X1 U4764 ( .A0(\reg_mem[12][4] ), .A1(\reg_mem[13][4] ), .S(net87388), 
        .Z(n3453) );
  CMXI2X1 U4765 ( .A0(\reg_mem[14][4] ), .A1(\reg_mem[15][4] ), .S(net87394), 
        .Z(n3452) );
  CMXI2X1 U4766 ( .A0(n3453), .A1(n3452), .S(n2176), .Z(n3454) );
  CMXI2X1 U4767 ( .A0(n3455), .A1(n3454), .S(net87247), .Z(n3456) );
  CMXI2X1 U4768 ( .A0(n3457), .A1(n3456), .S(net87522), .Z(n3471) );
  CMXI2X1 U4769 ( .A0(net79122), .A1(net79123), .S(n2182), .Z(n3461) );
  CMXI2X1 U4770 ( .A0(\reg_mem[20][4] ), .A1(\reg_mem[21][4] ), .S(net87387), 
        .Z(n3459) );
  CMXI2X1 U4771 ( .A0(\reg_mem[22][4] ), .A1(\reg_mem[23][4] ), .S(net87407), 
        .Z(n3458) );
  CMXI2X1 U4772 ( .A0(n3459), .A1(n3458), .S(n2183), .Z(n3460) );
  CMXI2X1 U4773 ( .A0(n3461), .A1(n3460), .S(net87247), .Z(n3469) );
  CMXI2X1 U4774 ( .A0(\reg_mem[24][4] ), .A1(\reg_mem[25][4] ), .S(net87411), 
        .Z(n3463) );
  CMXI2X1 U4775 ( .A0(\reg_mem[26][4] ), .A1(\reg_mem[27][4] ), .S(net87387), 
        .Z(n3462) );
  CMXI2X1 U4776 ( .A0(n3463), .A1(n3462), .S(n2197), .Z(n3467) );
  CMXI2X1 U4777 ( .A0(\reg_mem[28][4] ), .A1(\reg_mem[29][4] ), .S(net87412), 
        .Z(n3465) );
  CMXI2X1 U4778 ( .A0(\reg_mem[30][4] ), .A1(\reg_mem[31][4] ), .S(net87397), 
        .Z(n3464) );
  CMXI2X1 U4779 ( .A0(n3465), .A1(n3464), .S(n2190), .Z(n3466) );
  CMXI2X1 U4780 ( .A0(n3467), .A1(n3466), .S(net87272), .Z(n3468) );
  CMXI2X1 U4781 ( .A0(n3469), .A1(n3468), .S(net87523), .Z(n3470) );
  CIVX2 U4782 ( .A(alu_op_c[4]), .Z(n3472) );
  CIVX2 U4783 ( .A(N99), .Z(n3479) );
  CIVX2 U4784 ( .A(N67), .Z(n3474) );
  COND3X1 U4785 ( .A(n2115), .B(n3479), .C(n3478), .D(n3477), .Z(alu_op_c[3])
         );
  CND2IX1 U4786 ( .B(n2046), .A(n2146), .Z(n3485) );
  CND2IX1 U4787 ( .B(n3480), .A(n3741), .Z(n3483) );
  CMXI2X1 U4788 ( .A0(n3483), .A1(n3482), .S(prog_count_o[3]), .Z(n3484) );
  CMXI2X1 U4789 ( .A0(\reg_mem[0][3] ), .A1(\reg_mem[1][3] ), .S(net87407), 
        .Z(n3489) );
  CMXI2X1 U4790 ( .A0(n3489), .A1(n3488), .S(n2196), .Z(n3493) );
  CMXI2X1 U4791 ( .A0(\reg_mem[4][3] ), .A1(\reg_mem[5][3] ), .S(net87391), 
        .Z(n3491) );
  CMXI2X1 U4792 ( .A0(\reg_mem[6][3] ), .A1(\reg_mem[7][3] ), .S(net87387), 
        .Z(n3490) );
  CMXI2X1 U4793 ( .A0(n3491), .A1(n3490), .S(n2187), .Z(n3492) );
  CMXI2X1 U4794 ( .A0(\reg_mem[8][3] ), .A1(\reg_mem[9][3] ), .S(net87395), 
        .Z(n3495) );
  CMXI2X1 U4795 ( .A0(\reg_mem[10][3] ), .A1(\reg_mem[11][3] ), .S(net87407), 
        .Z(n3494) );
  CMXI2X1 U4796 ( .A0(n3495), .A1(n3494), .S(n2176), .Z(n3499) );
  CMXI2X1 U4797 ( .A0(\reg_mem[12][3] ), .A1(\reg_mem[13][3] ), .S(n2069), .Z(
        n3497) );
  CMXI2X1 U4798 ( .A0(\reg_mem[14][3] ), .A1(\reg_mem[15][3] ), .S(net87391), 
        .Z(n3496) );
  CMXI2X1 U4799 ( .A0(n3497), .A1(n3496), .S(n2177), .Z(n3498) );
  CMXI2X1 U4800 ( .A0(n3499), .A1(n3498), .S(net87268), .Z(n3500) );
  CMXI2X1 U4801 ( .A0(\reg_mem[16][3] ), .A1(\reg_mem[17][3] ), .S(net87398), 
        .Z(n3503) );
  CMXI2X1 U4802 ( .A0(\reg_mem[18][3] ), .A1(\reg_mem[19][3] ), .S(net87406), 
        .Z(n3502) );
  CMXI2X1 U4803 ( .A0(n3503), .A1(n3502), .S(n2181), .Z(n3507) );
  CMXI2X1 U4804 ( .A0(\reg_mem[20][3] ), .A1(\reg_mem[21][3] ), .S(net87399), 
        .Z(n3505) );
  CMXI2X1 U4805 ( .A0(\reg_mem[22][3] ), .A1(\reg_mem[23][3] ), .S(net87394), 
        .Z(n3504) );
  CMXI2X1 U4806 ( .A0(n3505), .A1(n3504), .S(n2182), .Z(n3506) );
  CMXI2X1 U4807 ( .A0(n3507), .A1(n3506), .S(n1480), .Z(n3515) );
  CMXI2X1 U4808 ( .A0(\reg_mem[24][3] ), .A1(\reg_mem[25][3] ), .S(net87401), 
        .Z(n3509) );
  CMXI2X1 U4809 ( .A0(\reg_mem[26][3] ), .A1(\reg_mem[27][3] ), .S(net87410), 
        .Z(n3508) );
  CMXI2X1 U4810 ( .A0(n3509), .A1(n3508), .S(n2196), .Z(n3513) );
  CMXI2X1 U4811 ( .A0(\reg_mem[28][3] ), .A1(\reg_mem[29][3] ), .S(net87392), 
        .Z(n3511) );
  CMXI2X1 U4812 ( .A0(\reg_mem[30][3] ), .A1(\reg_mem[31][3] ), .S(net87403), 
        .Z(n3510) );
  CMXI2X1 U4813 ( .A0(n3511), .A1(n3510), .S(n2166), .Z(n3512) );
  CMXI2X1 U4814 ( .A0(n3513), .A1(n3512), .S(net87271), .Z(n3514) );
  CMXI2X1 U4815 ( .A0(n3515), .A1(n3514), .S(net87856), .Z(n3516) );
  CIVX2 U4816 ( .A(alu_op_c[3]), .Z(n3518) );
  CANR2X1 U4817 ( .A(N171), .B(n3704), .C(N139), .D(n3701), .Z(n3521) );
  CMXI2X1 U4818 ( .A0(\reg_mem[0][2] ), .A1(\reg_mem[1][2] ), .S(net87400), 
        .Z(n3530) );
  CMXI2X1 U4819 ( .A0(\reg_mem[2][2] ), .A1(\reg_mem[3][2] ), .S(net87401), 
        .Z(n3529) );
  CMXI2X1 U4820 ( .A0(n3530), .A1(n3529), .S(n2195), .Z(n3534) );
  CMXI2X1 U4821 ( .A0(\reg_mem[4][2] ), .A1(\reg_mem[5][2] ), .S(net87389), 
        .Z(n3532) );
  CMXI2X1 U4822 ( .A0(\reg_mem[6][2] ), .A1(\reg_mem[7][2] ), .S(n1456), .Z(
        n3531) );
  CMXI2X1 U4823 ( .A0(n3532), .A1(n3531), .S(n2189), .Z(n3533) );
  CMXI2X1 U4824 ( .A0(n3534), .A1(n3533), .S(net87266), .Z(n3542) );
  CMXI2X1 U4825 ( .A0(\reg_mem[8][2] ), .A1(\reg_mem[9][2] ), .S(net87402), 
        .Z(n3536) );
  CMXI2X1 U4826 ( .A0(\reg_mem[10][2] ), .A1(\reg_mem[11][2] ), .S(net87389), 
        .Z(n3535) );
  CMXI2X1 U4827 ( .A0(n3536), .A1(n3535), .S(n2201), .Z(n3540) );
  CMXI2X1 U4828 ( .A0(\reg_mem[12][2] ), .A1(\reg_mem[13][2] ), .S(n2069), .Z(
        n3538) );
  CMXI2X1 U4829 ( .A0(\reg_mem[14][2] ), .A1(\reg_mem[15][2] ), .S(net87389), 
        .Z(n3537) );
  CMXI2X1 U4830 ( .A0(n3538), .A1(n3537), .S(n2201), .Z(n3539) );
  CMXI2X1 U4831 ( .A0(n3540), .A1(n3539), .S(net87275), .Z(n3541) );
  CMXI2X1 U4832 ( .A0(\reg_mem[20][2] ), .A1(\reg_mem[21][2] ), .S(net87393), 
        .Z(n3544) );
  CMXI2X1 U4833 ( .A0(\reg_mem[22][2] ), .A1(\reg_mem[23][2] ), .S(net87387), 
        .Z(n3543) );
  CMXI2X1 U4834 ( .A0(n3544), .A1(n3543), .S(n2181), .Z(n3545) );
  CMXI2X1 U4835 ( .A0(n3546), .A1(n3545), .S(n1385), .Z(n3554) );
  CMXI2X1 U4836 ( .A0(\reg_mem[24][2] ), .A1(\reg_mem[25][2] ), .S(net87398), 
        .Z(n3548) );
  CMXI2X1 U4837 ( .A0(\reg_mem[26][2] ), .A1(\reg_mem[27][2] ), .S(net87409), 
        .Z(n3547) );
  CMXI2X1 U4838 ( .A0(n3548), .A1(n3547), .S(n2195), .Z(n3552) );
  CMXI2X1 U4839 ( .A0(\reg_mem[28][2] ), .A1(\reg_mem[29][2] ), .S(net87387), 
        .Z(n3550) );
  CMXI2X1 U4840 ( .A0(\reg_mem[30][2] ), .A1(\reg_mem[31][2] ), .S(net87394), 
        .Z(n3549) );
  CMXI2X1 U4841 ( .A0(n3552), .A1(n3551), .S(n1480), .Z(n3553) );
  CMXI2X1 U4842 ( .A0(\reg_mem[0][1] ), .A1(\reg_mem[4][1] ), .S(net87242), 
        .Z(n3569) );
  CMXI2X1 U4843 ( .A0(\reg_mem[2][1] ), .A1(\reg_mem[6][1] ), .S(net87250), 
        .Z(n3568) );
  CMXI2X1 U4844 ( .A0(n3569), .A1(n3568), .S(n2193), .Z(n3573) );
  CMXI2X1 U4845 ( .A0(\reg_mem[1][1] ), .A1(\reg_mem[5][1] ), .S(net87250), 
        .Z(n3571) );
  CMXI2X1 U4846 ( .A0(\reg_mem[3][1] ), .A1(\reg_mem[7][1] ), .S(net87250), 
        .Z(n3570) );
  CMXI2X1 U4847 ( .A0(n3571), .A1(n3570), .S(n2189), .Z(n3572) );
  CMXI2X1 U4848 ( .A0(\reg_mem[10][1] ), .A1(\reg_mem[14][1] ), .S(net87250), 
        .Z(n3574) );
  CMXI2X1 U4849 ( .A0(\reg_mem[9][1] ), .A1(\reg_mem[13][1] ), .S(n1381), .Z(
        n3576) );
  CMXI2X1 U4850 ( .A0(\reg_mem[16][1] ), .A1(\reg_mem[17][1] ), .S(net87393), 
        .Z(n3582) );
  CMXI2X1 U4851 ( .A0(\reg_mem[18][1] ), .A1(\reg_mem[19][1] ), .S(net87395), 
        .Z(n3581) );
  CMXI2X1 U4852 ( .A0(n3582), .A1(n3581), .S(n2187), .Z(n3586) );
  CMXI2X1 U4853 ( .A0(\reg_mem[20][1] ), .A1(\reg_mem[21][1] ), .S(net87394), 
        .Z(n3584) );
  CMXI2X1 U4854 ( .A0(\reg_mem[22][1] ), .A1(\reg_mem[23][1] ), .S(net87397), 
        .Z(n3583) );
  CMXI2X1 U4855 ( .A0(n3586), .A1(n3585), .S(net87255), .Z(n3594) );
  CMXI2X1 U4856 ( .A0(\reg_mem[24][1] ), .A1(\reg_mem[25][1] ), .S(net87396), 
        .Z(n3588) );
  CMXI2X1 U4857 ( .A0(\reg_mem[26][1] ), .A1(\reg_mem[27][1] ), .S(net87398), 
        .Z(n3587) );
  CMXI2X1 U4858 ( .A0(n3588), .A1(n3587), .S(n2178), .Z(n3592) );
  CMXI2X1 U4859 ( .A0(\reg_mem[28][1] ), .A1(\reg_mem[29][1] ), .S(net87400), 
        .Z(n3590) );
  CMXI2X1 U4860 ( .A0(\reg_mem[30][1] ), .A1(\reg_mem[31][1] ), .S(net87401), 
        .Z(n3589) );
  CMXI2X1 U4861 ( .A0(n3590), .A1(n3589), .S(n2193), .Z(n3591) );
  CMXI2X1 U4862 ( .A0(n3592), .A1(n3591), .S(net87248), .Z(n3593) );
  CMXI2X1 U4863 ( .A0(n3594), .A1(n3593), .S(net87538), .Z(n3595) );
  CIVX2 U4864 ( .A(alu_op_c[1]), .Z(n3596) );
  CMXI2X1 U4865 ( .A0(\reg_mem[9][30] ), .A1(\reg_mem[25][30] ), .S(n2105), 
        .Z(n3598) );
  CMXI2X1 U4866 ( .A0(\reg_mem[11][30] ), .A1(\reg_mem[27][30] ), .S(n2090), 
        .Z(n3597) );
  CMXI2X1 U4867 ( .A0(n3598), .A1(n3597), .S(n2192), .Z(n3602) );
  CMXI2X1 U4868 ( .A0(\reg_mem[13][30] ), .A1(\reg_mem[29][30] ), .S(n1975), 
        .Z(n3600) );
  CMXI2X1 U4869 ( .A0(\reg_mem[2][30] ), .A1(\reg_mem[18][30] ), .S(n2104), 
        .Z(n3605) );
  CMXI2X1 U4870 ( .A0(n3606), .A1(n3605), .S(n2181), .Z(n3610) );
  CMXI2X1 U4871 ( .A0(\reg_mem[4][30] ), .A1(\reg_mem[20][30] ), .S(n2102), 
        .Z(n3608) );
  CMXI2X1 U4872 ( .A0(\reg_mem[6][30] ), .A1(\reg_mem[22][30] ), .S(n2092), 
        .Z(n3607) );
  CMXI2X1 U4873 ( .A0(n3608), .A1(n3607), .S(n2182), .Z(n3609) );
  CMXI2X1 U4874 ( .A0(n3610), .A1(n3609), .S(net87267), .Z(n3611) );
  CMXI2X1 U4875 ( .A0(\reg_mem[8][30] ), .A1(\reg_mem[24][30] ), .S(n2104), 
        .Z(n3617) );
  CMXI2X1 U4876 ( .A0(\reg_mem[10][30] ), .A1(\reg_mem[26][30] ), .S(n2093), 
        .Z(n3616) );
  CMXI2X1 U4877 ( .A0(\reg_mem[14][30] ), .A1(\reg_mem[30][30] ), .S(n2084), 
        .Z(n3618) );
  CMXI2X1 U4878 ( .A0(n3621), .A1(n3620), .S(net87271), .Z(n3622) );
  CND2IX1 U4879 ( .B(n3623), .A(n3622), .Z(n3633) );
  CMXI2X1 U4880 ( .A0(\reg_mem[1][30] ), .A1(\reg_mem[17][30] ), .S(n2101), 
        .Z(n3625) );
  CMXI2X1 U4881 ( .A0(\reg_mem[3][30] ), .A1(\reg_mem[19][30] ), .S(n2099), 
        .Z(n3624) );
  CMXI2X1 U4882 ( .A0(n3625), .A1(n3624), .S(n2190), .Z(n3629) );
  CMXI2X1 U4883 ( .A0(\reg_mem[7][30] ), .A1(\reg_mem[23][30] ), .S(n2087), 
        .Z(n3626) );
  CMXI2X1 U4884 ( .A0(n3629), .A1(n3628), .S(net87265), .Z(n3630) );
  CND2IX1 U4885 ( .B(n3631), .A(n3630), .Z(n3632) );
  CIVX2 U4886 ( .A(N126), .Z(n3634) );
  CND2IX1 U4887 ( .B(n3643), .A(n3642), .Z(alu_op_c[30]) );
  CND2IX1 U4888 ( .B(n3704), .A(n3690), .Z(n3645) );
  CMXI2X1 U4889 ( .A0(\reg_mem[5][31] ), .A1(\reg_mem[21][31] ), .S(n2092), 
        .Z(n3647) );
  CMXI2X1 U4890 ( .A0(n3647), .A1(n3646), .S(n2201), .Z(n3648) );
  CND2IX1 U4891 ( .B(n3649), .A(n3648), .Z(n3659) );
  CMXI2X1 U4892 ( .A0(\reg_mem[9][31] ), .A1(\reg_mem[25][31] ), .S(n2098), 
        .Z(n3651) );
  CND2IX1 U4893 ( .B(n3653), .A(n3652), .Z(n3658) );
  CMXI2X1 U4894 ( .A0(n3655), .A1(n3654), .S(n2166), .Z(n3656) );
  CANR1X1 U4895 ( .A(n2139), .B(n3656), .C(n1533), .Z(n3657) );
  CMXI2X1 U4896 ( .A0(\reg_mem[10][31] ), .A1(\reg_mem[26][31] ), .S(n1975), 
        .Z(n3660) );
  CND2IX1 U4897 ( .B(n3663), .A(n3662), .Z(n3674) );
  CMXI2X1 U4898 ( .A0(\reg_mem[12][31] ), .A1(\reg_mem[28][31] ), .S(n2082), 
        .Z(n3665) );
  CMXI2X1 U4899 ( .A0(\reg_mem[14][31] ), .A1(\reg_mem[30][31] ), .S(n2104), 
        .Z(n3664) );
  CMXI2X1 U4900 ( .A0(n3665), .A1(n3664), .S(n2192), .Z(n3666) );
  CND2IX1 U4901 ( .B(n3667), .A(n3666), .Z(n3673) );
  CMXI2X1 U4902 ( .A0(\reg_mem[1][31] ), .A1(\reg_mem[17][31] ), .S(n2088), 
        .Z(n3669) );
  CMXI2X1 U4903 ( .A0(n3669), .A1(n3668), .S(n2190), .Z(n3670) );
  CND2IX1 U4904 ( .B(n3671), .A(n3670), .Z(n3672) );
  CIVX2 U4905 ( .A(\reg_mem[0][31] ), .Z(n5160) );
  CIVX2 U4906 ( .A(\reg_mem[16][31] ), .Z(n5184) );
  CIVX2 U4907 ( .A(\reg_mem[2][31] ), .Z(n5162) );
  CIVX2 U4908 ( .A(\reg_mem[18][31] ), .Z(n5186) );
  CMXI2X1 U4909 ( .A0(n5162), .A1(n5186), .S(n2094), .Z(n3675) );
  CMXI2X1 U4910 ( .A0(n3676), .A1(n3675), .S(n2187), .Z(n3682) );
  CIVX2 U4911 ( .A(\reg_mem[4][31] ), .Z(n5166) );
  CIVX2 U4912 ( .A(\reg_mem[20][31] ), .Z(n5190) );
  CIVX2 U4913 ( .A(\reg_mem[6][31] ), .Z(n5168) );
  CIVX2 U4914 ( .A(\reg_mem[22][31] ), .Z(n5192) );
  CMXI2X1 U4915 ( .A0(n5168), .A1(n5192), .S(n2083), .Z(n3677) );
  CMXI2X1 U4916 ( .A0(n3678), .A1(n3677), .S(n2186), .Z(n3680) );
  COND2X2 U4917 ( .A(n3682), .B(n3681), .C(n3680), .D(n3679), .Z(n3683) );
  CIVX2 U4918 ( .A(N72), .Z(n3698) );
  CANR2X1 U4919 ( .A(N145), .B(n3701), .C(n2157), .D(n3700), .Z(n3702) );
  CIVX2 U4920 ( .A(n3702), .Z(n3703) );
  CMXI2X1 U4921 ( .A0(\reg_mem[6][8] ), .A1(\reg_mem[7][8] ), .S(net87404), 
        .Z(n3710) );
  CMXI2X1 U4922 ( .A0(n3712), .A1(n3711), .S(net87260), .Z(n3720) );
  CMXI2X1 U4923 ( .A0(\reg_mem[8][8] ), .A1(\reg_mem[9][8] ), .S(net87404), 
        .Z(n3714) );
  CMXI2X1 U4924 ( .A0(\reg_mem[10][8] ), .A1(\reg_mem[11][8] ), .S(net87388), 
        .Z(n3713) );
  CMXI2X1 U4925 ( .A0(n3714), .A1(n3713), .S(n2192), .Z(n3718) );
  CMXI2X1 U4926 ( .A0(\reg_mem[12][8] ), .A1(\reg_mem[13][8] ), .S(net87408), 
        .Z(n3716) );
  CMXI2X1 U4927 ( .A0(\reg_mem[14][8] ), .A1(\reg_mem[15][8] ), .S(net87406), 
        .Z(n3715) );
  CMXI2X1 U4928 ( .A0(n3716), .A1(n3715), .S(n2176), .Z(n3717) );
  CMXI2X1 U4929 ( .A0(n3718), .A1(n3717), .S(n1385), .Z(n3719) );
  CMXI2X1 U4930 ( .A0(\reg_mem[16][8] ), .A1(\reg_mem[17][8] ), .S(net87400), 
        .Z(n3722) );
  CMXI2X1 U4931 ( .A0(\reg_mem[18][8] ), .A1(\reg_mem[19][8] ), .S(net87403), 
        .Z(n3721) );
  CMXI2X1 U4932 ( .A0(n3722), .A1(n3721), .S(n2165), .Z(n3726) );
  CMXI2X1 U4933 ( .A0(\reg_mem[20][8] ), .A1(\reg_mem[21][8] ), .S(n1456), .Z(
        n3724) );
  CMXI2X1 U4934 ( .A0(\reg_mem[22][8] ), .A1(\reg_mem[23][8] ), .S(n2069), .Z(
        n3723) );
  CMXI2X1 U4935 ( .A0(n3724), .A1(n3723), .S(n2166), .Z(n3725) );
  CMXI2X1 U4936 ( .A0(n3726), .A1(n3725), .S(n1480), .Z(n3734) );
  CMXI2X1 U4937 ( .A0(\reg_mem[24][8] ), .A1(\reg_mem[25][8] ), .S(net87405), 
        .Z(n3728) );
  CMXI2X1 U4938 ( .A0(\reg_mem[26][8] ), .A1(\reg_mem[27][8] ), .S(net87408), 
        .Z(n3727) );
  CMXI2X1 U4939 ( .A0(n3728), .A1(n3727), .S(n2166), .Z(n3732) );
  CMXI2X1 U4940 ( .A0(\reg_mem[28][8] ), .A1(\reg_mem[29][8] ), .S(n2069), .Z(
        n3730) );
  CMXI2X1 U4941 ( .A0(\reg_mem[30][8] ), .A1(\reg_mem[31][8] ), .S(net87401), 
        .Z(n3729) );
  CMXI2X1 U4942 ( .A0(n3730), .A1(n3729), .S(n2191), .Z(n3731) );
  CMXI2X1 U4943 ( .A0(n3732), .A1(n3731), .S(net87252), .Z(n3733) );
  CMXI2X1 U4944 ( .A0(n3734), .A1(n3733), .S(n1532), .Z(n3735) );
  CIVX2 U4945 ( .A(alu_op_c[8]), .Z(n3737) );
  CANR2X1 U4946 ( .A(alu_op_c[7]), .B(n3750), .C(regA[7]), .D(n3739), .Z(n3749) );
  CIVX2 U4947 ( .A(prog_count_o[6]), .Z(n3740) );
  CND2IX1 U4948 ( .B(n3740), .A(n2155), .Z(n3745) );
  CND2IX1 U4949 ( .B(prog_count_o[6]), .A(n3741), .Z(n3743) );
  CMXI2X1 U4950 ( .A0(n3745), .A1(n3744), .S(prog_count_o[7]), .Z(n3746) );
  CIVX2 U4951 ( .A(n5235), .Z(n5237) );
  CIVX2 U4952 ( .A(n5262), .Z(n5217) );
  CIVX2 U4953 ( .A(n5261), .Z(n5218) );
  CIVX2 U4954 ( .A(n5260), .Z(n5219) );
  CIVX2 U4955 ( .A(n5259), .Z(n5220) );
  CIVX2 U4956 ( .A(n5258), .Z(n5221) );
  CIVX2 U4957 ( .A(n5257), .Z(n5222) );
  CIVX2 U4958 ( .A(n5256), .Z(n5223) );
  CIVX2 U4959 ( .A(n5255), .Z(n5224) );
  CIVX2 U4960 ( .A(n5254), .Z(n5225) );
  CIVX2 U4961 ( .A(n5253), .Z(n5226) );
  CIVX2 U4962 ( .A(n5252), .Z(n5227) );
  CMXI2X1 U4963 ( .A0(n3758), .A1(n3757), .S(net87640), .Z(n3764) );
  CIVX2 U4964 ( .A(\reg_mem[6][0] ), .Z(n3760) );
  CIVX2 U4965 ( .A(\reg_mem[7][0] ), .Z(n3759) );
  CMXI2X1 U4966 ( .A0(n3760), .A1(n3759), .S(net87804), .Z(n3761) );
  CMXI2X1 U4967 ( .A0(n3762), .A1(n3761), .S(net87623), .Z(n3763) );
  CMXI2X1 U4968 ( .A0(n3764), .A1(n3763), .S(net87727), .Z(n3774) );
  CMXI2X1 U4969 ( .A0(n3766), .A1(n3765), .S(net87636), .Z(n3772) );
  CIVX2 U4970 ( .A(\reg_mem[14][0] ), .Z(n3768) );
  CIVX2 U4971 ( .A(\reg_mem[15][0] ), .Z(n3767) );
  CMXI2X1 U4972 ( .A0(n3768), .A1(n3767), .S(net87794), .Z(n3769) );
  CMXI2X1 U4973 ( .A0(n3770), .A1(n3769), .S(net87627), .Z(n3771) );
  CMXI2X1 U4974 ( .A0(n3772), .A1(n3771), .S(net87724), .Z(n3773) );
  CMXI2X1 U4975 ( .A0(n3774), .A1(n3773), .S(net82859), .Z(n3800) );
  CMXI2X1 U4976 ( .A0(n3776), .A1(n3775), .S(net87629), .Z(n3782) );
  CIVX2 U4977 ( .A(\reg_mem[22][0] ), .Z(n3778) );
  CIVX2 U4978 ( .A(\reg_mem[23][0] ), .Z(n3777) );
  CMXI2X1 U4979 ( .A0(n3778), .A1(n3777), .S(net87793), .Z(n3779) );
  CIVX2 U4980 ( .A(\reg_mem[24][0] ), .Z(n3784) );
  CIVX2 U4981 ( .A(\reg_mem[25][0] ), .Z(n3783) );
  CMXI2X1 U4982 ( .A0(n3784), .A1(n3783), .S(net87795), .Z(n3788) );
  CIVX2 U4983 ( .A(\reg_mem[26][0] ), .Z(n3786) );
  CIVX2 U4984 ( .A(\reg_mem[27][0] ), .Z(n3785) );
  CMXI2X1 U4985 ( .A0(n3786), .A1(n3785), .S(net87798), .Z(n3787) );
  CMXI2X1 U4986 ( .A0(n3788), .A1(n3787), .S(net87635), .Z(n3796) );
  CIVX2 U4987 ( .A(\reg_mem[28][0] ), .Z(n3790) );
  CMXI2X1 U4988 ( .A0(n3790), .A1(n3789), .S(net87807), .Z(n3794) );
  CIVX2 U4989 ( .A(\reg_mem[30][0] ), .Z(n3792) );
  CIVX2 U4990 ( .A(\reg_mem[31][0] ), .Z(n3791) );
  CMXI2X1 U4991 ( .A0(n3792), .A1(n3791), .S(net87794), .Z(n3793) );
  CMXI2X1 U4992 ( .A0(n3794), .A1(n3793), .S(net87625), .Z(n3795) );
  CMXI2X1 U4993 ( .A0(n3796), .A1(n3795), .S(net87717), .Z(n3797) );
  CMXI2X1 U4994 ( .A0(n3802), .A1(n3801), .S(net87632), .Z(n3808) );
  CIVX2 U4995 ( .A(\reg_mem[6][1] ), .Z(n3804) );
  CIVX2 U4996 ( .A(\reg_mem[7][1] ), .Z(n3803) );
  CMXI2X1 U4997 ( .A0(n3804), .A1(n3803), .S(net87800), .Z(n3805) );
  CMXI2X1 U4998 ( .A0(n3806), .A1(n3805), .S(net87639), .Z(n3807) );
  CMXI2X1 U4999 ( .A0(n3808), .A1(n3807), .S(net87716), .Z(n3818) );
  CMXI2X1 U5000 ( .A0(n3810), .A1(n3809), .S(net87632), .Z(n3816) );
  CIVX2 U5001 ( .A(\reg_mem[14][1] ), .Z(n3812) );
  CIVX2 U5002 ( .A(\reg_mem[15][1] ), .Z(n3811) );
  CMXI2X1 U5003 ( .A0(n3812), .A1(n3811), .S(net87791), .Z(n3813) );
  CMXI2X1 U5004 ( .A0(n3814), .A1(n3813), .S(net87634), .Z(n3815) );
  CMXI2X1 U5005 ( .A0(n3816), .A1(n3815), .S(net87727), .Z(n3817) );
  CMXI2X1 U5006 ( .A0(n3818), .A1(n3817), .S(net82859), .Z(n3844) );
  CMXI2X1 U5007 ( .A0(n3820), .A1(n3819), .S(net87635), .Z(n3826) );
  CIVX2 U5008 ( .A(\reg_mem[22][1] ), .Z(n3822) );
  CIVX2 U5009 ( .A(\reg_mem[23][1] ), .Z(n3821) );
  CMXI2X1 U5010 ( .A0(n3822), .A1(n3821), .S(net87800), .Z(n3823) );
  CMXI2X1 U5011 ( .A0(n3824), .A1(n3823), .S(net87637), .Z(n3825) );
  CMXI2X1 U5012 ( .A0(n3826), .A1(n3825), .S(net87708), .Z(n3842) );
  CIVX2 U5013 ( .A(\reg_mem[24][1] ), .Z(n3828) );
  CIVX2 U5014 ( .A(\reg_mem[25][1] ), .Z(n3827) );
  CMXI2X1 U5015 ( .A0(n3828), .A1(n3827), .S(net87799), .Z(n3832) );
  CIVX2 U5016 ( .A(\reg_mem[26][1] ), .Z(n3830) );
  CIVX2 U5017 ( .A(\reg_mem[27][1] ), .Z(n3829) );
  CMXI2X1 U5018 ( .A0(n3832), .A1(n3831), .S(net87636), .Z(n3840) );
  CIVX2 U5019 ( .A(\reg_mem[28][1] ), .Z(n3834) );
  CMXI2X1 U5020 ( .A0(n3834), .A1(n3833), .S(net87794), .Z(n3838) );
  CIVX2 U5021 ( .A(\reg_mem[30][1] ), .Z(n3836) );
  CIVX2 U5022 ( .A(\reg_mem[31][1] ), .Z(n3835) );
  CMXI2X1 U5023 ( .A0(n3836), .A1(n3835), .S(net87809), .Z(n3837) );
  CMXI2X1 U5024 ( .A0(n3838), .A1(n3837), .S(net87638), .Z(n3839) );
  CMXI2X1 U5025 ( .A0(n3840), .A1(n3839), .S(net87719), .Z(n3841) );
  CMXI2X1 U5026 ( .A0(n3842), .A1(n3841), .S(net82859), .Z(n3843) );
  CMXI2X1 U5027 ( .A0(n3844), .A1(n3843), .S(net86657), .Z(N231) );
  CMXI2X1 U5028 ( .A0(n3846), .A1(n3845), .S(net87635), .Z(n3852) );
  CIVX2 U5029 ( .A(\reg_mem[6][2] ), .Z(n3848) );
  CIVX2 U5030 ( .A(\reg_mem[7][2] ), .Z(n3847) );
  CMXI2X1 U5031 ( .A0(n3848), .A1(n3847), .S(net87791), .Z(n3849) );
  CMXI2X1 U5032 ( .A0(n3850), .A1(n3849), .S(net87630), .Z(n3851) );
  CMXI2X1 U5033 ( .A0(n3852), .A1(n3851), .S(net87725), .Z(n3862) );
  CIVX2 U5034 ( .A(\reg_mem[14][2] ), .Z(n3856) );
  CIVX2 U5035 ( .A(\reg_mem[15][2] ), .Z(n3855) );
  CMXI2X1 U5036 ( .A0(n3856), .A1(n3855), .S(net87797), .Z(n3857) );
  CMXI2X1 U5037 ( .A0(n3860), .A1(n3859), .S(net87728), .Z(n3861) );
  CIVX2 U5038 ( .A(\reg_mem[22][2] ), .Z(net78621) );
  CIVX2 U5039 ( .A(\reg_mem[23][2] ), .Z(net78622) );
  CIVX2 U5040 ( .A(\reg_mem[24][2] ), .Z(n3864) );
  CIVX2 U5041 ( .A(\reg_mem[25][2] ), .Z(n3863) );
  CMXI2X1 U5042 ( .A0(n3864), .A1(n3863), .S(net87806), .Z(n3868) );
  CIVX2 U5043 ( .A(\reg_mem[26][2] ), .Z(n3866) );
  CIVX2 U5044 ( .A(\reg_mem[27][2] ), .Z(n3865) );
  CMXI2X1 U5045 ( .A0(n3866), .A1(n3865), .S(net87795), .Z(n3867) );
  CMXI2X1 U5046 ( .A0(n3868), .A1(n3867), .S(net87632), .Z(n3876) );
  CIVX2 U5047 ( .A(\reg_mem[28][2] ), .Z(n3870) );
  CMXI2X1 U5048 ( .A0(n3870), .A1(n3869), .S(net87795), .Z(n3874) );
  CIVX2 U5049 ( .A(\reg_mem[30][2] ), .Z(n3872) );
  CIVX2 U5050 ( .A(\reg_mem[31][2] ), .Z(n3871) );
  CMXI2X1 U5051 ( .A0(n3872), .A1(n3871), .S(net87806), .Z(n3873) );
  CMXI2X1 U5052 ( .A0(n3874), .A1(n3873), .S(net87624), .Z(n3875) );
  CMXI2X1 U5053 ( .A0(n3876), .A1(n3875), .S(net87706), .Z(net78602) );
  CMXI2X1 U5054 ( .A0(n3878), .A1(n3877), .S(net87639), .Z(n3884) );
  CIVX2 U5055 ( .A(\reg_mem[6][3] ), .Z(n3880) );
  CIVX2 U5056 ( .A(\reg_mem[7][3] ), .Z(n3879) );
  CMXI2X1 U5057 ( .A0(n3880), .A1(n3879), .S(net87806), .Z(n3881) );
  CMXI2X1 U5058 ( .A0(n3882), .A1(n3881), .S(net87642), .Z(n3883) );
  CMXI2X1 U5059 ( .A0(n3884), .A1(n3883), .S(net87724), .Z(n3894) );
  CMXI2X1 U5060 ( .A0(n3886), .A1(n3885), .S(net87634), .Z(n3892) );
  CIVX2 U5061 ( .A(\reg_mem[14][3] ), .Z(n3888) );
  CIVX2 U5062 ( .A(\reg_mem[15][3] ), .Z(n3887) );
  CMXI2X1 U5063 ( .A0(n3888), .A1(n3887), .S(net87806), .Z(n3889) );
  CMXI2X1 U5064 ( .A0(n3890), .A1(n3889), .S(net87626), .Z(n3891) );
  CMXI2X1 U5065 ( .A0(n3892), .A1(n3891), .S(net87727), .Z(n3893) );
  CMXI2X1 U5066 ( .A0(n3894), .A1(n3893), .S(net82859), .Z(n3920) );
  CIVX2 U5067 ( .A(\reg_mem[22][3] ), .Z(n3898) );
  CIVX2 U5068 ( .A(\reg_mem[23][3] ), .Z(n3897) );
  CMXI2X1 U5069 ( .A0(n3898), .A1(n3897), .S(net87804), .Z(n3899) );
  CMXI2X1 U5070 ( .A0(n3902), .A1(n3901), .S(net87705), .Z(n3918) );
  CIVX2 U5071 ( .A(\reg_mem[24][3] ), .Z(n3904) );
  CIVX2 U5072 ( .A(\reg_mem[25][3] ), .Z(n3903) );
  CMXI2X1 U5073 ( .A0(n3904), .A1(n3903), .S(net87794), .Z(n3908) );
  CIVX2 U5074 ( .A(\reg_mem[26][3] ), .Z(n3906) );
  CIVX2 U5075 ( .A(\reg_mem[27][3] ), .Z(n3905) );
  CMXI2X1 U5076 ( .A0(n3906), .A1(n3905), .S(net87804), .Z(n3907) );
  CMXI2X1 U5077 ( .A0(n3908), .A1(n3907), .S(net87625), .Z(n3916) );
  CIVX2 U5078 ( .A(\reg_mem[28][3] ), .Z(n3910) );
  CMXI2X1 U5079 ( .A0(n3910), .A1(n3909), .S(net87793), .Z(n3914) );
  CIVX2 U5080 ( .A(\reg_mem[30][3] ), .Z(n3912) );
  CIVX2 U5081 ( .A(\reg_mem[31][3] ), .Z(n3911) );
  CMXI2X1 U5082 ( .A0(n3912), .A1(n3911), .S(net87799), .Z(n3913) );
  CMXI2X1 U5083 ( .A0(n3914), .A1(n3913), .S(net87624), .Z(n3915) );
  CMXI2X1 U5084 ( .A0(n3916), .A1(n3915), .S(net87705), .Z(n3917) );
  CIVX2 U5085 ( .A(\reg_mem[6][4] ), .Z(n3924) );
  CIVX2 U5086 ( .A(\reg_mem[7][4] ), .Z(n3923) );
  CMXI2X1 U5087 ( .A0(n3924), .A1(n3923), .S(net87800), .Z(n3925) );
  CMXI2X1 U5088 ( .A0(n3926), .A1(n3925), .S(net87634), .Z(n3927) );
  CMXI2X1 U5089 ( .A0(n3928), .A1(n3927), .S(net87728), .Z(n3938) );
  CMXI2X1 U5090 ( .A0(n3930), .A1(n3929), .S(net87631), .Z(n3936) );
  CIVX2 U5091 ( .A(\reg_mem[14][4] ), .Z(n3932) );
  CIVX2 U5092 ( .A(\reg_mem[15][4] ), .Z(n3931) );
  CMXI2X1 U5093 ( .A0(n3932), .A1(n3931), .S(net87804), .Z(n3933) );
  CMXI2X1 U5094 ( .A0(n3934), .A1(n3933), .S(net87631), .Z(n3935) );
  CMXI2X1 U5095 ( .A0(n3936), .A1(n3935), .S(net87705), .Z(n3937) );
  CMXI2X1 U5096 ( .A0(n3938), .A1(n3937), .S(net82859), .Z(net78475) );
  CIVX2 U5097 ( .A(\reg_mem[22][4] ), .Z(net78497) );
  CIVX2 U5098 ( .A(\reg_mem[23][4] ), .Z(net78498) );
  CIVX2 U5099 ( .A(\reg_mem[24][4] ), .Z(n3940) );
  CIVX2 U5100 ( .A(\reg_mem[25][4] ), .Z(n3939) );
  CMXI2X1 U5101 ( .A0(n3940), .A1(n3939), .S(net87807), .Z(n3944) );
  CIVX2 U5102 ( .A(\reg_mem[26][4] ), .Z(n3942) );
  CIVX2 U5103 ( .A(\reg_mem[27][4] ), .Z(n3941) );
  CMXI2X1 U5104 ( .A0(n3942), .A1(n3941), .S(net87794), .Z(n3943) );
  CMXI2X1 U5105 ( .A0(n3944), .A1(n3943), .S(net87633), .Z(n3952) );
  CIVX2 U5106 ( .A(\reg_mem[28][4] ), .Z(n3946) );
  CMXI2X1 U5107 ( .A0(n3946), .A1(n3945), .S(net87797), .Z(n3950) );
  CIVX2 U5108 ( .A(\reg_mem[30][4] ), .Z(n3948) );
  CIVX2 U5109 ( .A(\reg_mem[31][4] ), .Z(n3947) );
  CMXI2X1 U5110 ( .A0(n3948), .A1(n3947), .S(net87809), .Z(n3949) );
  CMXI2X1 U5111 ( .A0(n3950), .A1(n3949), .S(net87640), .Z(n3951) );
  CMXI2X1 U5112 ( .A0(n3952), .A1(n3951), .S(net87709), .Z(net78478) );
  CMXI2X1 U5113 ( .A0(n3954), .A1(n3953), .S(net87629), .Z(n3960) );
  CIVX2 U5114 ( .A(\reg_mem[6][5] ), .Z(n3956) );
  CIVX2 U5115 ( .A(\reg_mem[7][5] ), .Z(n3955) );
  CMXI2X1 U5116 ( .A0(n3956), .A1(n3955), .S(net87803), .Z(n3957) );
  CMXI2X1 U5117 ( .A0(n3958), .A1(n3957), .S(net87630), .Z(n3959) );
  CMXI2X1 U5118 ( .A0(n3962), .A1(n3961), .S(net87630), .Z(n3968) );
  CIVX2 U5119 ( .A(\reg_mem[14][5] ), .Z(n3964) );
  CIVX2 U5120 ( .A(\reg_mem[15][5] ), .Z(n3963) );
  CMXI2X1 U5121 ( .A0(n3964), .A1(n3963), .S(net87793), .Z(n3965) );
  CMXI2X1 U5122 ( .A0(n3972), .A1(n3971), .S(net87629), .Z(n3978) );
  CIVX2 U5123 ( .A(\reg_mem[22][5] ), .Z(n3974) );
  CIVX2 U5124 ( .A(\reg_mem[23][5] ), .Z(n3973) );
  CMXI2X1 U5125 ( .A0(n3974), .A1(n3973), .S(net87791), .Z(n3975) );
  CMXI2X1 U5126 ( .A0(n3978), .A1(n3977), .S(net87704), .Z(n3994) );
  CIVX2 U5127 ( .A(\reg_mem[24][5] ), .Z(n3980) );
  CIVX2 U5128 ( .A(\reg_mem[25][5] ), .Z(n3979) );
  CMXI2X1 U5129 ( .A0(n3980), .A1(n3979), .S(net87804), .Z(n3984) );
  CIVX2 U5130 ( .A(\reg_mem[26][5] ), .Z(n3982) );
  CIVX2 U5131 ( .A(\reg_mem[27][5] ), .Z(n3981) );
  CMXI2X1 U5132 ( .A0(n3984), .A1(n3983), .S(net87631), .Z(n3992) );
  CIVX2 U5133 ( .A(\reg_mem[28][5] ), .Z(n3986) );
  CMXI2X1 U5134 ( .A0(n3986), .A1(n3985), .S(net87807), .Z(n3990) );
  CIVX2 U5135 ( .A(\reg_mem[30][5] ), .Z(n3988) );
  CMXI2X1 U5136 ( .A0(n3988), .A1(n3987), .S(net87795), .Z(n3989) );
  CMXI2X1 U5137 ( .A0(n3990), .A1(n3989), .S(net87628), .Z(n3991) );
  CMXI2X1 U5138 ( .A0(n3992), .A1(n3991), .S(net87730), .Z(n3993) );
  CMXI2X1 U5139 ( .A0(n3994), .A1(n3993), .S(net82859), .Z(n3995) );
  CMXI2X1 U5140 ( .A0(n3998), .A1(n3997), .S(net87631), .Z(n4004) );
  CIVX2 U5141 ( .A(\reg_mem[6][6] ), .Z(n4000) );
  CIVX2 U5142 ( .A(\reg_mem[7][6] ), .Z(n3999) );
  CMXI2X1 U5143 ( .A0(n4004), .A1(n4003), .S(net87705), .Z(n4014) );
  CIVX2 U5144 ( .A(\reg_mem[14][6] ), .Z(n4008) );
  CIVX2 U5145 ( .A(\reg_mem[15][6] ), .Z(n4007) );
  CMXI2X1 U5146 ( .A0(n4012), .A1(n4011), .S(net87724), .Z(n4013) );
  CIVX2 U5147 ( .A(\reg_mem[22][6] ), .Z(n4018) );
  CIVX2 U5148 ( .A(\reg_mem[23][6] ), .Z(n4017) );
  CMXI2X1 U5149 ( .A0(n4020), .A1(n4019), .S(net87629), .Z(n4021) );
  CMXI2X1 U5150 ( .A0(n4022), .A1(n4021), .S(net87730), .Z(n4038) );
  CIVX2 U5151 ( .A(\reg_mem[24][6] ), .Z(n4024) );
  CIVX2 U5152 ( .A(\reg_mem[25][6] ), .Z(n4023) );
  CIVX2 U5153 ( .A(\reg_mem[26][6] ), .Z(n4026) );
  CIVX2 U5154 ( .A(\reg_mem[27][6] ), .Z(n4025) );
  CMXI2X1 U5155 ( .A0(n4026), .A1(n4025), .S(net87802), .Z(n4027) );
  CMXI2X1 U5156 ( .A0(n4028), .A1(n4027), .S(net87625), .Z(n4036) );
  CIVX2 U5157 ( .A(\reg_mem[28][6] ), .Z(n4030) );
  CMXI2X1 U5158 ( .A0(n4030), .A1(n4029), .S(net87802), .Z(n4034) );
  CIVX2 U5159 ( .A(\reg_mem[30][6] ), .Z(n4032) );
  CIVX2 U5160 ( .A(\reg_mem[31][6] ), .Z(n4031) );
  CMXI2X1 U5161 ( .A0(n4032), .A1(n4031), .S(net87803), .Z(n4033) );
  CMXI2X1 U5162 ( .A0(n4034), .A1(n4033), .S(net87633), .Z(n4035) );
  CMXI2X1 U5163 ( .A0(n4036), .A1(n4035), .S(net87724), .Z(n4037) );
  CMXI2X1 U5164 ( .A0(n4038), .A1(n4037), .S(net82861), .Z(n4039) );
  CMXI2X1 U5165 ( .A0(n4042), .A1(n4041), .S(net87636), .Z(n4048) );
  CIVX2 U5166 ( .A(\reg_mem[6][7] ), .Z(n4044) );
  CIVX2 U5167 ( .A(\reg_mem[7][7] ), .Z(n4043) );
  CMXI2X1 U5168 ( .A0(n4044), .A1(n4043), .S(net87806), .Z(n4045) );
  CMXI2X1 U5169 ( .A0(n4046), .A1(n4045), .S(net87631), .Z(n4047) );
  CMXI2X1 U5170 ( .A0(n4048), .A1(n4047), .S(net87720), .Z(n4058) );
  CMXI2X1 U5171 ( .A0(n4050), .A1(n4049), .S(net87638), .Z(n4056) );
  CIVX2 U5172 ( .A(\reg_mem[14][7] ), .Z(n4052) );
  CIVX2 U5173 ( .A(\reg_mem[15][7] ), .Z(n4051) );
  CMXI2X1 U5174 ( .A0(n4052), .A1(n4051), .S(net87798), .Z(n4053) );
  CMXI2X1 U5175 ( .A0(n4054), .A1(n4053), .S(net87640), .Z(n4055) );
  CMXI2X1 U5176 ( .A0(n4056), .A1(n4055), .S(net87725), .Z(n4057) );
  CMXI2X1 U5177 ( .A0(n4058), .A1(n4057), .S(net82861), .Z(n4084) );
  CMXI2X1 U5178 ( .A0(n4060), .A1(n4059), .S(net87639), .Z(n4066) );
  CIVX2 U5179 ( .A(\reg_mem[22][7] ), .Z(n4062) );
  CIVX2 U5180 ( .A(\reg_mem[23][7] ), .Z(n4061) );
  CMXI2X1 U5181 ( .A0(n4062), .A1(n4061), .S(net87802), .Z(n4063) );
  CMXI2X1 U5182 ( .A0(n4066), .A1(n4065), .S(net87728), .Z(n4082) );
  CIVX2 U5183 ( .A(\reg_mem[24][7] ), .Z(n4068) );
  CIVX2 U5184 ( .A(\reg_mem[25][7] ), .Z(n4067) );
  CMXI2X1 U5185 ( .A0(n4068), .A1(n4067), .S(net87799), .Z(n4072) );
  CIVX2 U5186 ( .A(\reg_mem[26][7] ), .Z(n4070) );
  CIVX2 U5187 ( .A(\reg_mem[27][7] ), .Z(n4069) );
  CMXI2X1 U5188 ( .A0(n4070), .A1(n4069), .S(net87799), .Z(n4071) );
  CIVX2 U5189 ( .A(\reg_mem[28][7] ), .Z(n4074) );
  CMXI2X1 U5190 ( .A0(n4074), .A1(n4073), .S(net87793), .Z(n4078) );
  CIVX2 U5191 ( .A(\reg_mem[30][7] ), .Z(n4076) );
  CMXI2X1 U5192 ( .A0(n4076), .A1(n4075), .S(net87803), .Z(n4077) );
  CMXI2X1 U5193 ( .A0(n4080), .A1(n4079), .S(net87716), .Z(n4081) );
  CIVX2 U5194 ( .A(\reg_mem[0][8] ), .Z(n4086) );
  CIVX2 U5195 ( .A(\reg_mem[1][8] ), .Z(n4085) );
  CIVX2 U5196 ( .A(\reg_mem[6][8] ), .Z(n4090) );
  CIVX2 U5197 ( .A(\reg_mem[7][8] ), .Z(n4089) );
  CMXI2X1 U5198 ( .A0(n4090), .A1(n4089), .S(net87807), .Z(n4091) );
  CMXI2X1 U5199 ( .A0(n4094), .A1(n4093), .S(net87719), .Z(n4104) );
  CIVX2 U5200 ( .A(\reg_mem[14][8] ), .Z(n4098) );
  CIVX2 U5201 ( .A(\reg_mem[15][8] ), .Z(n4097) );
  CMXI2X1 U5202 ( .A0(n4098), .A1(n4097), .S(net87806), .Z(n4099) );
  CMXI2X1 U5203 ( .A0(n4102), .A1(n4101), .S(net87724), .Z(n4103) );
  CMXI2X1 U5204 ( .A0(n4104), .A1(n4103), .S(net82861), .Z(n4130) );
  CMXI2X1 U5205 ( .A0(n4106), .A1(n4105), .S(net87632), .Z(n4112) );
  CIVX2 U5206 ( .A(\reg_mem[22][8] ), .Z(n4108) );
  CIVX2 U5207 ( .A(\reg_mem[23][8] ), .Z(n4107) );
  CMXI2X1 U5208 ( .A0(n4108), .A1(n4107), .S(net87798), .Z(n4109) );
  CMXI2X1 U5209 ( .A0(n4110), .A1(n4109), .S(net87628), .Z(n4111) );
  CMXI2X1 U5210 ( .A0(n4112), .A1(n4111), .S(net87730), .Z(n4128) );
  CIVX2 U5211 ( .A(\reg_mem[24][8] ), .Z(n4114) );
  CIVX2 U5212 ( .A(\reg_mem[25][8] ), .Z(n4113) );
  CMXI2X1 U5213 ( .A0(n4114), .A1(n4113), .S(net87807), .Z(n4118) );
  CIVX2 U5214 ( .A(\reg_mem[26][8] ), .Z(n4116) );
  CIVX2 U5215 ( .A(\reg_mem[27][8] ), .Z(n4115) );
  CMXI2X1 U5216 ( .A0(n4116), .A1(n4115), .S(net87803), .Z(n4117) );
  CMXI2X1 U5217 ( .A0(n4118), .A1(n4117), .S(net87636), .Z(n4126) );
  CIVX2 U5218 ( .A(\reg_mem[28][8] ), .Z(n4120) );
  CMXI2X1 U5219 ( .A0(n4120), .A1(n4119), .S(net87797), .Z(n4124) );
  CIVX2 U5220 ( .A(\reg_mem[30][8] ), .Z(n4122) );
  CIVX2 U5221 ( .A(\reg_mem[31][8] ), .Z(n4121) );
  CMXI2X1 U5222 ( .A0(n4122), .A1(n4121), .S(net87794), .Z(n4123) );
  CMXI2X1 U5223 ( .A0(n4124), .A1(n4123), .S(net87626), .Z(n4125) );
  CMXI2X1 U5224 ( .A0(n4126), .A1(n4125), .S(net87710), .Z(n4127) );
  CMXI2X1 U5225 ( .A0(n4128), .A1(n4127), .S(net82861), .Z(n4129) );
  CIVX2 U5226 ( .A(\reg_mem[6][9] ), .Z(n4134) );
  CIVX2 U5227 ( .A(\reg_mem[7][9] ), .Z(n4133) );
  CMXI2X1 U5228 ( .A0(n4134), .A1(n4133), .S(net87798), .Z(n4135) );
  CMXI2X1 U5229 ( .A0(n4136), .A1(n4135), .S(net87626), .Z(n4137) );
  CMXI2X1 U5230 ( .A0(n4140), .A1(n4139), .S(net87624), .Z(n4146) );
  CIVX2 U5231 ( .A(\reg_mem[14][9] ), .Z(n4142) );
  CIVX2 U5232 ( .A(\reg_mem[15][9] ), .Z(n4141) );
  CMXI2X1 U5233 ( .A0(n4142), .A1(n4141), .S(net87791), .Z(n4143) );
  CMXI2X1 U5234 ( .A0(n4146), .A1(n4145), .S(net87715), .Z(n4147) );
  CMXI2X1 U5235 ( .A0(n4148), .A1(n4147), .S(net82861), .Z(n4174) );
  CIVX2 U5236 ( .A(\reg_mem[22][9] ), .Z(n4152) );
  CIVX2 U5237 ( .A(\reg_mem[23][9] ), .Z(n4151) );
  CMXI2X1 U5238 ( .A0(n4152), .A1(n4151), .S(net87791), .Z(n4153) );
  CMXI2X1 U5239 ( .A0(n4154), .A1(n4153), .S(net87629), .Z(n4155) );
  CIVX2 U5240 ( .A(\reg_mem[24][9] ), .Z(n4158) );
  CIVX2 U5241 ( .A(\reg_mem[25][9] ), .Z(n4157) );
  CMXI2X1 U5242 ( .A0(n4158), .A1(n4157), .S(net87802), .Z(n4162) );
  CIVX2 U5243 ( .A(\reg_mem[26][9] ), .Z(n4160) );
  CIVX2 U5244 ( .A(\reg_mem[27][9] ), .Z(n4159) );
  CMXI2X1 U5245 ( .A0(n4160), .A1(n4159), .S(net87807), .Z(n4161) );
  CIVX2 U5246 ( .A(\reg_mem[28][9] ), .Z(n4164) );
  CMXI2X1 U5247 ( .A0(n4164), .A1(n4163), .S(net87797), .Z(n4168) );
  CIVX2 U5248 ( .A(\reg_mem[30][9] ), .Z(n4166) );
  CIVX2 U5249 ( .A(\reg_mem[31][9] ), .Z(n4165) );
  CMXI2X1 U5250 ( .A0(n4166), .A1(n4165), .S(net87800), .Z(n4167) );
  CMXI2X1 U5251 ( .A0(n4168), .A1(n4167), .S(net87630), .Z(n4169) );
  CMXI2X1 U5252 ( .A0(n4170), .A1(n4169), .S(net87704), .Z(n4171) );
  CMXI2X1 U5253 ( .A0(n4176), .A1(n4175), .S(net87631), .Z(n4182) );
  CIVX2 U5254 ( .A(\reg_mem[6][10] ), .Z(n4178) );
  CIVX2 U5255 ( .A(\reg_mem[7][10] ), .Z(n4177) );
  CMXI2X1 U5256 ( .A0(n4178), .A1(n4177), .S(net87800), .Z(n4179) );
  CMXI2X1 U5257 ( .A0(n4180), .A1(n4179), .S(net87640), .Z(n4181) );
  CMXI2X1 U5258 ( .A0(n4184), .A1(n4183), .S(net87642), .Z(n4190) );
  CIVX2 U5259 ( .A(\reg_mem[14][10] ), .Z(n4186) );
  CIVX2 U5260 ( .A(\reg_mem[15][10] ), .Z(n4185) );
  CMXI2X1 U5261 ( .A0(n4186), .A1(n4185), .S(net87795), .Z(n4187) );
  CMXI2X1 U5262 ( .A0(n4188), .A1(n4187), .S(net87638), .Z(n4189) );
  CMXI2X1 U5263 ( .A0(n4190), .A1(n4189), .S(net87723), .Z(n4191) );
  CMXI2X1 U5264 ( .A0(n4192), .A1(n4191), .S(net82861), .Z(n4218) );
  CMXI2X1 U5265 ( .A0(n4194), .A1(n4193), .S(net87627), .Z(n4200) );
  CIVX2 U5266 ( .A(\reg_mem[22][10] ), .Z(n4196) );
  CIVX2 U5267 ( .A(\reg_mem[23][10] ), .Z(n4195) );
  CMXI2X1 U5268 ( .A0(n4196), .A1(n4195), .S(net87791), .Z(n4197) );
  CMXI2X1 U5269 ( .A0(n4198), .A1(n4197), .S(net87625), .Z(n4199) );
  CIVX2 U5270 ( .A(\reg_mem[24][10] ), .Z(n4202) );
  CIVX2 U5271 ( .A(\reg_mem[25][10] ), .Z(n4201) );
  CMXI2X1 U5272 ( .A0(n4202), .A1(n4201), .S(net87802), .Z(n4206) );
  CIVX2 U5273 ( .A(\reg_mem[26][10] ), .Z(n4204) );
  CIVX2 U5274 ( .A(\reg_mem[27][10] ), .Z(n4203) );
  CMXI2X1 U5275 ( .A0(n4204), .A1(n4203), .S(net87793), .Z(n4205) );
  CMXI2X1 U5276 ( .A0(n4206), .A1(n4205), .S(net87624), .Z(n4214) );
  CIVX2 U5277 ( .A(\reg_mem[28][10] ), .Z(n4208) );
  CMXI2X1 U5278 ( .A0(n4208), .A1(n4207), .S(net87794), .Z(n4212) );
  CIVX2 U5279 ( .A(\reg_mem[30][10] ), .Z(n4210) );
  CIVX2 U5280 ( .A(\reg_mem[31][10] ), .Z(n4209) );
  CMXI2X1 U5281 ( .A0(n4212), .A1(n4211), .S(net87623), .Z(n4213) );
  CMXI2X1 U5282 ( .A0(n4214), .A1(n4213), .S(net87709), .Z(n4215) );
  CMXI2X1 U5283 ( .A0(n4216), .A1(n4215), .S(net82861), .Z(n4217) );
  CIVX2 U5284 ( .A(\reg_mem[14][11] ), .Z(n4222) );
  CIVX2 U5285 ( .A(\reg_mem[15][11] ), .Z(n4221) );
  CMXI2X1 U5286 ( .A0(n4226), .A1(n4225), .S(net87722), .Z(net78074) );
  CMXI2X1 U5287 ( .A0(n4228), .A1(n4227), .S(net87626), .Z(n4234) );
  CIVX2 U5288 ( .A(\reg_mem[22][11] ), .Z(n4230) );
  CIVX2 U5289 ( .A(\reg_mem[23][11] ), .Z(n4229) );
  CMXI2X1 U5290 ( .A0(n4230), .A1(n4229), .S(net87809), .Z(n4231) );
  CMXI2X1 U5291 ( .A0(n4232), .A1(n4231), .S(net87624), .Z(n4233) );
  CMXI2X1 U5292 ( .A0(n4234), .A1(n4233), .S(net87728), .Z(n4250) );
  CIVX2 U5293 ( .A(\reg_mem[24][11] ), .Z(n4236) );
  CIVX2 U5294 ( .A(\reg_mem[25][11] ), .Z(n4235) );
  CMXI2X1 U5295 ( .A0(n4236), .A1(n4235), .S(net87797), .Z(n4240) );
  CIVX2 U5296 ( .A(\reg_mem[26][11] ), .Z(n4238) );
  CIVX2 U5297 ( .A(\reg_mem[27][11] ), .Z(n4237) );
  CMXI2X1 U5298 ( .A0(n4238), .A1(n4237), .S(net87809), .Z(n4239) );
  CMXI2X1 U5299 ( .A0(n4240), .A1(n4239), .S(net87636), .Z(n4248) );
  CIVX2 U5300 ( .A(\reg_mem[28][11] ), .Z(n4242) );
  CMXI2X1 U5301 ( .A0(n4242), .A1(n4241), .S(net87809), .Z(n4246) );
  CIVX2 U5302 ( .A(\reg_mem[30][11] ), .Z(n4244) );
  CIVX2 U5303 ( .A(\reg_mem[31][11] ), .Z(n4243) );
  CMXI2X1 U5304 ( .A0(n4244), .A1(n4243), .S(net87800), .Z(n4245) );
  CMXI2X1 U5305 ( .A0(n4246), .A1(n4245), .S(net87642), .Z(n4247) );
  CMXI2X1 U5306 ( .A0(n4248), .A1(n4247), .S(net87708), .Z(n4249) );
  CMXI2X1 U5307 ( .A0(n4250), .A1(n4249), .S(net82861), .Z(net78042) );
  CIVX2 U5308 ( .A(\reg_mem[6][12] ), .Z(n4254) );
  CIVX2 U5309 ( .A(\reg_mem[7][12] ), .Z(n4253) );
  CMXI2X1 U5310 ( .A0(n4254), .A1(n4253), .S(net87803), .Z(n4255) );
  CMXI2X1 U5311 ( .A0(n4258), .A1(n4257), .S(net87716), .Z(n4268) );
  CIVX2 U5312 ( .A(\reg_mem[14][12] ), .Z(n4262) );
  CIVX2 U5313 ( .A(\reg_mem[15][12] ), .Z(n4261) );
  CMXI2X1 U5314 ( .A0(n4262), .A1(n4261), .S(net87794), .Z(n4263) );
  CMXI2X1 U5315 ( .A0(n4264), .A1(n4263), .S(net87642), .Z(n4265) );
  CMXI2X1 U5316 ( .A0(n4266), .A1(n4265), .S(net87722), .Z(n4267) );
  CMXI2X1 U5317 ( .A0(n4270), .A1(n4269), .S(net87638), .Z(n4276) );
  CIVX2 U5318 ( .A(\reg_mem[22][12] ), .Z(n4272) );
  CIVX2 U5319 ( .A(\reg_mem[23][12] ), .Z(n4271) );
  CMXI2X1 U5320 ( .A0(n4272), .A1(n4271), .S(net87803), .Z(n4273) );
  CMXI2X1 U5321 ( .A0(n4274), .A1(n4273), .S(net87640), .Z(n4275) );
  CIVX2 U5322 ( .A(\reg_mem[24][12] ), .Z(n4278) );
  CIVX2 U5323 ( .A(\reg_mem[25][12] ), .Z(n4277) );
  CMXI2X1 U5324 ( .A0(n4278), .A1(n4277), .S(net87806), .Z(n4282) );
  CIVX2 U5325 ( .A(\reg_mem[26][12] ), .Z(n4280) );
  CIVX2 U5326 ( .A(\reg_mem[27][12] ), .Z(n4279) );
  CMXI2X1 U5327 ( .A0(n4280), .A1(n4279), .S(net87798), .Z(n4281) );
  CIVX2 U5328 ( .A(\reg_mem[28][12] ), .Z(n4284) );
  CMXI2X1 U5329 ( .A0(n4284), .A1(n4283), .S(net87794), .Z(n4288) );
  CIVX2 U5330 ( .A(\reg_mem[30][12] ), .Z(n4286) );
  CIVX2 U5331 ( .A(\reg_mem[31][12] ), .Z(n4285) );
  CMXI2X1 U5332 ( .A0(n4286), .A1(n4285), .S(net87804), .Z(n4287) );
  CMXI2X1 U5333 ( .A0(n4290), .A1(n4289), .S(net87725), .Z(n4291) );
  CMXI2X1 U5334 ( .A0(n4296), .A1(n4295), .S(net87628), .Z(n4302) );
  CIVX2 U5335 ( .A(\reg_mem[14][13] ), .Z(n4298) );
  CIVX2 U5336 ( .A(\reg_mem[15][13] ), .Z(n4297) );
  CMXI2X1 U5337 ( .A0(n4298), .A1(n4297), .S(net87799), .Z(n4299) );
  CMXI2X1 U5338 ( .A0(n4300), .A1(n4299), .S(net87624), .Z(n4301) );
  CMXI2X1 U5339 ( .A0(n4304), .A1(n4303), .S(net87625), .Z(n4310) );
  CIVX2 U5340 ( .A(\reg_mem[22][13] ), .Z(n4306) );
  CIVX2 U5341 ( .A(\reg_mem[23][13] ), .Z(n4305) );
  CMXI2X1 U5342 ( .A0(n4306), .A1(n4305), .S(net87802), .Z(n4307) );
  CMXI2X1 U5343 ( .A0(n4308), .A1(n4307), .S(net87623), .Z(n4309) );
  CMXI2X1 U5344 ( .A0(n4310), .A1(n4309), .S(net87724), .Z(n4326) );
  CIVX2 U5345 ( .A(\reg_mem[24][13] ), .Z(n4312) );
  CIVX2 U5346 ( .A(\reg_mem[25][13] ), .Z(n4311) );
  CMXI2X1 U5347 ( .A0(n4312), .A1(n4311), .S(net87797), .Z(n4316) );
  CIVX2 U5348 ( .A(\reg_mem[26][13] ), .Z(n4314) );
  CIVX2 U5349 ( .A(\reg_mem[27][13] ), .Z(n4313) );
  CMXI2X1 U5350 ( .A0(n4314), .A1(n4313), .S(net87800), .Z(n4315) );
  CMXI2X1 U5351 ( .A0(n4316), .A1(n4315), .S(net87634), .Z(n4324) );
  CIVX2 U5352 ( .A(\reg_mem[28][13] ), .Z(n4318) );
  CMXI2X1 U5353 ( .A0(n4318), .A1(n4317), .S(net87791), .Z(n4322) );
  CIVX2 U5354 ( .A(\reg_mem[30][13] ), .Z(n4320) );
  CIVX2 U5355 ( .A(\reg_mem[31][13] ), .Z(n4319) );
  CMXI2X1 U5356 ( .A0(n4320), .A1(n4319), .S(net87795), .Z(n4321) );
  CMXI2X1 U5357 ( .A0(n4324), .A1(n4323), .S(net87706), .Z(n4325) );
  CMXI2X1 U5358 ( .A0(n4328), .A1(n4327), .S(net87631), .Z(n4334) );
  CIVX2 U5359 ( .A(\reg_mem[6][14] ), .Z(n4330) );
  CIVX2 U5360 ( .A(\reg_mem[7][14] ), .Z(n4329) );
  CMXI2X1 U5361 ( .A0(n4330), .A1(n4329), .S(net87798), .Z(n4331) );
  CMXI2X1 U5362 ( .A0(n4332), .A1(n4331), .S(net87638), .Z(n4333) );
  CMXI2X1 U5363 ( .A0(n4334), .A1(n4333), .S(net87715), .Z(n4344) );
  CIVX2 U5364 ( .A(\reg_mem[14][14] ), .Z(n4338) );
  CIVX2 U5365 ( .A(\reg_mem[15][14] ), .Z(n4337) );
  CMXI2X1 U5366 ( .A0(n4338), .A1(n4337), .S(net87791), .Z(n4339) );
  CMXI2X1 U5367 ( .A0(n4340), .A1(n4339), .S(net87633), .Z(n4341) );
  CMXI2X1 U5368 ( .A0(n4344), .A1(n4343), .S(net82863), .Z(n4370) );
  CMXI2X1 U5369 ( .A0(n4346), .A1(n4345), .S(net87628), .Z(n4352) );
  CIVX2 U5370 ( .A(\reg_mem[22][14] ), .Z(n4348) );
  CIVX2 U5371 ( .A(\reg_mem[23][14] ), .Z(n4347) );
  CMXI2X1 U5372 ( .A0(n4348), .A1(n4347), .S(net87799), .Z(n4349) );
  CMXI2X1 U5373 ( .A0(n4350), .A1(n4349), .S(net87636), .Z(n4351) );
  CMXI2X1 U5374 ( .A0(n4352), .A1(n4351), .S(net87710), .Z(n4368) );
  CIVX2 U5375 ( .A(\reg_mem[24][14] ), .Z(n4354) );
  CIVX2 U5376 ( .A(\reg_mem[25][14] ), .Z(n4353) );
  CMXI2X1 U5377 ( .A0(n4354), .A1(n4353), .S(net87807), .Z(n4358) );
  CIVX2 U5378 ( .A(\reg_mem[26][14] ), .Z(n4356) );
  CIVX2 U5379 ( .A(\reg_mem[27][14] ), .Z(n4355) );
  CMXI2X1 U5380 ( .A0(n4356), .A1(n4355), .S(net87803), .Z(n4357) );
  CMXI2X1 U5381 ( .A0(n4358), .A1(n4357), .S(net87625), .Z(n4366) );
  CIVX2 U5382 ( .A(\reg_mem[28][14] ), .Z(n4360) );
  CMXI2X1 U5383 ( .A0(n4360), .A1(n4359), .S(net87803), .Z(n4364) );
  CIVX2 U5384 ( .A(\reg_mem[30][14] ), .Z(n4362) );
  CIVX2 U5385 ( .A(\reg_mem[31][14] ), .Z(n4361) );
  CMXI2X1 U5386 ( .A0(n4362), .A1(n4361), .S(net87809), .Z(n4363) );
  CMXI2X1 U5387 ( .A0(n4364), .A1(n4363), .S(net87625), .Z(n4365) );
  CMXI2X1 U5388 ( .A0(n4366), .A1(n4365), .S(net87718), .Z(n4367) );
  CMXI2X1 U5389 ( .A0(n4368), .A1(n4367), .S(net82863), .Z(n4369) );
  CIVX2 U5390 ( .A(\reg_mem[0][15] ), .Z(n4372) );
  CMXI2X1 U5391 ( .A0(n4372), .A1(n4371), .S(net87800), .Z(n4376) );
  CIVX2 U5392 ( .A(\reg_mem[2][15] ), .Z(n4374) );
  CMXI2X1 U5393 ( .A0(n4374), .A1(n4373), .S(net87799), .Z(n4375) );
  CMXI2X1 U5394 ( .A0(n4376), .A1(n4375), .S(net87636), .Z(n4384) );
  CIVX2 U5395 ( .A(\reg_mem[4][15] ), .Z(n4378) );
  CMXI2X1 U5396 ( .A0(n4378), .A1(n4377), .S(net87793), .Z(n4382) );
  CIVX2 U5397 ( .A(\reg_mem[6][15] ), .Z(n4380) );
  CMXI2X1 U5398 ( .A0(n4380), .A1(n4379), .S(net87807), .Z(n4381) );
  CMXI2X1 U5399 ( .A0(n4382), .A1(n4381), .S(net87635), .Z(n4383) );
  CMXI2X1 U5400 ( .A0(n4384), .A1(n4383), .S(net87714), .Z(n4400) );
  CMXI2X1 U5401 ( .A0(n4386), .A1(n4385), .S(net87807), .Z(n4390) );
  CMXI2X1 U5402 ( .A0(n4388), .A1(n4387), .S(net87802), .Z(n4389) );
  CMXI2X1 U5403 ( .A0(n4390), .A1(n4389), .S(net87627), .Z(n4398) );
  CMXI2X1 U5404 ( .A0(n4392), .A1(n4391), .S(net87794), .Z(n4396) );
  CMXI2X1 U5405 ( .A0(n4394), .A1(n4393), .S(net87807), .Z(n4395) );
  CMXI2X1 U5406 ( .A0(n4396), .A1(n4395), .S(net87640), .Z(n4397) );
  CMXI2X1 U5407 ( .A0(n4398), .A1(n4397), .S(net87722), .Z(n4399) );
  CMXI2X1 U5408 ( .A0(n4400), .A1(n4399), .S(net82863), .Z(n4432) );
  CIVX2 U5409 ( .A(\reg_mem[16][15] ), .Z(n4402) );
  CIVX2 U5410 ( .A(\reg_mem[18][15] ), .Z(n4404) );
  CMXI2X1 U5411 ( .A0(n4404), .A1(n4403), .S(net87795), .Z(n4405) );
  CIVX2 U5412 ( .A(\reg_mem[20][15] ), .Z(n4408) );
  CMXI2X1 U5413 ( .A0(n4408), .A1(n4407), .S(net87804), .Z(n4412) );
  CIVX2 U5414 ( .A(\reg_mem[22][15] ), .Z(n4410) );
  CMXI2X1 U5415 ( .A0(n4410), .A1(n4409), .S(net87794), .Z(n4411) );
  CMXI2X1 U5416 ( .A0(n4412), .A1(n4411), .S(net87639), .Z(n4413) );
  CMXI2X1 U5417 ( .A0(n4414), .A1(n4413), .S(net87725), .Z(n4430) );
  CMXI2X1 U5418 ( .A0(n4418), .A1(n4417), .S(net87791), .Z(n4419) );
  CMXI2X1 U5419 ( .A0(n4420), .A1(n4419), .S(net87626), .Z(n4428) );
  CMXI2X1 U5420 ( .A0(n4422), .A1(n4421), .S(net87804), .Z(n4426) );
  CMXI2X1 U5421 ( .A0(n4424), .A1(n4423), .S(net87794), .Z(n4425) );
  CMXI2X1 U5422 ( .A0(n4426), .A1(n4425), .S(net87637), .Z(n4427) );
  CMXI2X1 U5423 ( .A0(n4428), .A1(n4427), .S(net87705), .Z(n4429) );
  CMXI2X1 U5424 ( .A0(n4430), .A1(n4429), .S(net82863), .Z(n4431) );
  CMXI2X1 U5425 ( .A0(n4432), .A1(n4431), .S(net86657), .Z(N217) );
  CIVX2 U5426 ( .A(\reg_mem[6][16] ), .Z(n4434) );
  CIVX2 U5427 ( .A(\reg_mem[7][16] ), .Z(n4433) );
  CMXI2X1 U5428 ( .A0(n4434), .A1(n4433), .S(net87800), .Z(n4435) );
  CMXI2X1 U5429 ( .A0(n4436), .A1(n4435), .S(net87633), .Z(n4437) );
  CMXI2X1 U5430 ( .A0(n4438), .A1(n4437), .S(net87727), .Z(n4448) );
  CMXI2X1 U5431 ( .A0(n4440), .A1(n4439), .S(net87630), .Z(n4446) );
  CIVX2 U5432 ( .A(\reg_mem[14][16] ), .Z(n4442) );
  CIVX2 U5433 ( .A(\reg_mem[15][16] ), .Z(n4441) );
  CMXI2X1 U5434 ( .A0(n4442), .A1(n4441), .S(net87804), .Z(n4443) );
  CMXI2X1 U5435 ( .A0(n4444), .A1(n4443), .S(net87630), .Z(n4445) );
  CMXI2X1 U5436 ( .A0(n4446), .A1(n4445), .S(net87730), .Z(n4447) );
  CMXI2X1 U5437 ( .A0(n4448), .A1(n4447), .S(net82863), .Z(n4474) );
  CMXI2X1 U5438 ( .A0(n4450), .A1(n4449), .S(net87632), .Z(n4456) );
  CIVX2 U5439 ( .A(\reg_mem[22][16] ), .Z(n4452) );
  CIVX2 U5440 ( .A(\reg_mem[23][16] ), .Z(n4451) );
  CMXI2X1 U5441 ( .A0(n4452), .A1(n4451), .S(net87803), .Z(n4453) );
  CMXI2X1 U5442 ( .A0(n4454), .A1(n4453), .S(net87633), .Z(n4455) );
  CIVX2 U5443 ( .A(\reg_mem[24][16] ), .Z(n4458) );
  CIVX2 U5444 ( .A(\reg_mem[25][16] ), .Z(n4457) );
  CMXI2X1 U5445 ( .A0(n4458), .A1(n4457), .S(net87806), .Z(n4462) );
  CIVX2 U5446 ( .A(\reg_mem[26][16] ), .Z(n4460) );
  CIVX2 U5447 ( .A(\reg_mem[27][16] ), .Z(n4459) );
  CMXI2X1 U5448 ( .A0(n4460), .A1(n4459), .S(net87800), .Z(n4461) );
  CMXI2X1 U5449 ( .A0(n4462), .A1(n4461), .S(net87635), .Z(n4470) );
  CIVX2 U5450 ( .A(\reg_mem[28][16] ), .Z(n4464) );
  CIVX2 U5451 ( .A(\reg_mem[29][16] ), .Z(n4463) );
  CMXI2X1 U5452 ( .A0(n4464), .A1(n4463), .S(net87791), .Z(n4468) );
  CIVX2 U5453 ( .A(\reg_mem[30][16] ), .Z(n4466) );
  CIVX2 U5454 ( .A(\reg_mem[31][16] ), .Z(n4465) );
  CMXI2X1 U5455 ( .A0(n4466), .A1(n4465), .S(net87807), .Z(n4467) );
  CMXI2X1 U5456 ( .A0(n4468), .A1(n4467), .S(net87638), .Z(n4469) );
  CMXI2X1 U5457 ( .A0(n4470), .A1(n4469), .S(net87708), .Z(n4471) );
  CMXI2X1 U5458 ( .A0(n4472), .A1(n4471), .S(net82863), .Z(n4473) );
  CMXI2X1 U5459 ( .A0(n4476), .A1(n4475), .S(net87633), .Z(n4482) );
  CIVX2 U5460 ( .A(\reg_mem[6][17] ), .Z(n4478) );
  CIVX2 U5461 ( .A(\reg_mem[7][17] ), .Z(n4477) );
  CMXI2X1 U5462 ( .A0(n4478), .A1(n4477), .S(net87806), .Z(n4479) );
  CMXI2X1 U5463 ( .A0(n4480), .A1(n4479), .S(net87640), .Z(n4481) );
  CIVX2 U5464 ( .A(\reg_mem[14][17] ), .Z(n4486) );
  CIVX2 U5465 ( .A(\reg_mem[15][17] ), .Z(n4485) );
  CMXI2X1 U5466 ( .A0(n4486), .A1(n4485), .S(net87799), .Z(n4487) );
  CMXI2X1 U5467 ( .A0(n4488), .A1(n4487), .S(net87625), .Z(n4489) );
  CMXI2X1 U5468 ( .A0(n4490), .A1(n4489), .S(net87718), .Z(n4491) );
  CIVX2 U5469 ( .A(\reg_mem[22][17] ), .Z(n4496) );
  CIVX2 U5470 ( .A(\reg_mem[23][17] ), .Z(n4495) );
  CMXI2X1 U5471 ( .A0(n4496), .A1(n4495), .S(net87809), .Z(n4497) );
  CMXI2X1 U5472 ( .A0(n4498), .A1(n4497), .S(net87626), .Z(n4499) );
  CIVX2 U5473 ( .A(\reg_mem[24][17] ), .Z(n4502) );
  CIVX2 U5474 ( .A(\reg_mem[25][17] ), .Z(n4501) );
  CMXI2X1 U5475 ( .A0(n4502), .A1(n4501), .S(net87800), .Z(n4506) );
  CIVX2 U5476 ( .A(\reg_mem[26][17] ), .Z(n4504) );
  CIVX2 U5477 ( .A(\reg_mem[27][17] ), .Z(n4503) );
  CMXI2X1 U5478 ( .A0(n4504), .A1(n4503), .S(net87800), .Z(n4505) );
  CMXI2X1 U5479 ( .A0(n4506), .A1(n4505), .S(net87633), .Z(n4514) );
  CIVX2 U5480 ( .A(\reg_mem[28][17] ), .Z(n4508) );
  CIVX2 U5481 ( .A(\reg_mem[29][17] ), .Z(n4507) );
  CMXI2X1 U5482 ( .A0(n4508), .A1(n4507), .S(net87800), .Z(n4512) );
  CIVX2 U5483 ( .A(\reg_mem[30][17] ), .Z(n4510) );
  CIVX2 U5484 ( .A(\reg_mem[31][17] ), .Z(n4509) );
  CMXI2X1 U5485 ( .A0(n4510), .A1(n4509), .S(net87794), .Z(n4511) );
  CMXI2X1 U5486 ( .A0(n4512), .A1(n4511), .S(net87640), .Z(n4513) );
  CMXI2X1 U5487 ( .A0(n4514), .A1(n4513), .S(net87704), .Z(n4515) );
  CIVX2 U5488 ( .A(\reg_mem[6][18] ), .Z(n4522) );
  CIVX2 U5489 ( .A(\reg_mem[7][18] ), .Z(n4521) );
  CMXI2X1 U5490 ( .A0(n4522), .A1(n4521), .S(net87797), .Z(n4523) );
  CMXI2X1 U5491 ( .A0(n4524), .A1(n4523), .S(net87627), .Z(n4525) );
  CMXI2X1 U5492 ( .A0(n4526), .A1(n4525), .S(net87714), .Z(n4536) );
  CIVX2 U5493 ( .A(\reg_mem[14][18] ), .Z(n4530) );
  CIVX2 U5494 ( .A(\reg_mem[15][18] ), .Z(n4529) );
  CMXI2X1 U5495 ( .A0(n4530), .A1(n4529), .S(net87797), .Z(n4531) );
  CMXI2X1 U5496 ( .A0(n4532), .A1(n4531), .S(net87629), .Z(n4533) );
  CMXI2X1 U5497 ( .A0(n4534), .A1(n4533), .S(net87716), .Z(n4535) );
  CIVX2 U5498 ( .A(\reg_mem[22][18] ), .Z(n4540) );
  CIVX2 U5499 ( .A(\reg_mem[23][18] ), .Z(n4539) );
  CMXI2X1 U5500 ( .A0(n4540), .A1(n4539), .S(net87791), .Z(n4541) );
  CMXI2X1 U5501 ( .A0(n4542), .A1(n4541), .S(net87633), .Z(n4543) );
  CMXI2X1 U5502 ( .A0(n4544), .A1(n4543), .S(net87709), .Z(n4560) );
  CIVX2 U5503 ( .A(\reg_mem[24][18] ), .Z(n4546) );
  CIVX2 U5504 ( .A(\reg_mem[25][18] ), .Z(n4545) );
  CMXI2X1 U5505 ( .A0(n4546), .A1(n4545), .S(net87800), .Z(n4550) );
  CIVX2 U5506 ( .A(\reg_mem[26][18] ), .Z(n4548) );
  CIVX2 U5507 ( .A(\reg_mem[27][18] ), .Z(n4547) );
  CMXI2X1 U5508 ( .A0(n4548), .A1(n4547), .S(net87791), .Z(n4549) );
  CMXI2X1 U5509 ( .A0(n4550), .A1(n4549), .S(net87628), .Z(n4558) );
  CIVX2 U5510 ( .A(\reg_mem[28][18] ), .Z(n4552) );
  CIVX2 U5511 ( .A(\reg_mem[29][18] ), .Z(n4551) );
  CMXI2X1 U5512 ( .A0(n4552), .A1(n4551), .S(net87798), .Z(n4556) );
  CIVX2 U5513 ( .A(\reg_mem[30][18] ), .Z(n4554) );
  CIVX2 U5514 ( .A(\reg_mem[31][18] ), .Z(n4553) );
  CMXI2X1 U5515 ( .A0(n4554), .A1(n4553), .S(net87793), .Z(n4555) );
  CMXI2X1 U5516 ( .A0(n4556), .A1(n4555), .S(net87634), .Z(n4557) );
  CMXI2X1 U5517 ( .A0(n4558), .A1(n4557), .S(net87717), .Z(n4559) );
  CMXI2X1 U5518 ( .A0(n4564), .A1(n4563), .S(net87624), .Z(n4570) );
  CIVX2 U5519 ( .A(\reg_mem[6][19] ), .Z(n4566) );
  CIVX2 U5520 ( .A(\reg_mem[7][19] ), .Z(n4565) );
  CMXI2X1 U5521 ( .A0(n4566), .A1(n4565), .S(net87807), .Z(n4567) );
  CIVX2 U5522 ( .A(\reg_mem[14][19] ), .Z(n4572) );
  CIVX2 U5523 ( .A(\reg_mem[15][19] ), .Z(n4571) );
  CMXI2X1 U5524 ( .A0(n4572), .A1(n4571), .S(net87807), .Z(n4573) );
  CMXI2X1 U5525 ( .A0(n4574), .A1(n4573), .S(net87634), .Z(n4575) );
  CMXI2X1 U5526 ( .A0(n4576), .A1(n4575), .S(net87720), .Z(n4577) );
  CMXI2X1 U5527 ( .A0(n4578), .A1(n4577), .S(net82865), .Z(n4602) );
  CIVX2 U5528 ( .A(\reg_mem[22][19] ), .Z(n4580) );
  CIVX2 U5529 ( .A(\reg_mem[23][19] ), .Z(n4579) );
  CMXI2X1 U5530 ( .A0(n4580), .A1(n4579), .S(net87793), .Z(n4581) );
  CMXI2X1 U5531 ( .A0(n4584), .A1(n4583), .S(net87723), .Z(n4600) );
  CIVX2 U5532 ( .A(\reg_mem[24][19] ), .Z(n4586) );
  CIVX2 U5533 ( .A(\reg_mem[25][19] ), .Z(n4585) );
  CMXI2X1 U5534 ( .A0(n4586), .A1(n4585), .S(net87799), .Z(n4590) );
  CIVX2 U5535 ( .A(\reg_mem[26][19] ), .Z(n4588) );
  CIVX2 U5536 ( .A(\reg_mem[27][19] ), .Z(n4587) );
  CMXI2X1 U5537 ( .A0(n4588), .A1(n4587), .S(net87794), .Z(n4589) );
  CMXI2X1 U5538 ( .A0(n4590), .A1(n4589), .S(net87632), .Z(n4598) );
  CIVX2 U5539 ( .A(\reg_mem[28][19] ), .Z(n4592) );
  CIVX2 U5540 ( .A(\reg_mem[29][19] ), .Z(n4591) );
  CMXI2X1 U5541 ( .A0(n4592), .A1(n4591), .S(net87797), .Z(n4596) );
  CIVX2 U5542 ( .A(\reg_mem[30][19] ), .Z(n4594) );
  CIVX2 U5543 ( .A(\reg_mem[31][19] ), .Z(n4593) );
  CMXI2X1 U5544 ( .A0(n4594), .A1(n4593), .S(net87791), .Z(n4595) );
  CMXI2X1 U5545 ( .A0(n4596), .A1(n4595), .S(net87629), .Z(n4597) );
  CMXI2X1 U5546 ( .A0(n4598), .A1(n4597), .S(net87704), .Z(n4599) );
  CMXI2X1 U5547 ( .A0(n4604), .A1(n4603), .S(net87632), .Z(n4610) );
  CIVX2 U5548 ( .A(\reg_mem[6][20] ), .Z(n4606) );
  CIVX2 U5549 ( .A(\reg_mem[7][20] ), .Z(n4605) );
  CMXI2X1 U5550 ( .A0(n4606), .A1(n4605), .S(net87802), .Z(n4607) );
  CMXI2X1 U5551 ( .A0(n4608), .A1(n4607), .S(net87639), .Z(n4609) );
  CIVX2 U5552 ( .A(\reg_mem[14][20] ), .Z(n4614) );
  CIVX2 U5553 ( .A(\reg_mem[15][20] ), .Z(n4613) );
  CMXI2X1 U5554 ( .A0(n4614), .A1(n4613), .S(net87804), .Z(n4615) );
  CMXI2X1 U5555 ( .A0(n4618), .A1(n4617), .S(net87719), .Z(n4619) );
  CMXI2X1 U5556 ( .A0(n4622), .A1(n4621), .S(net87642), .Z(n4628) );
  CIVX2 U5557 ( .A(\reg_mem[22][20] ), .Z(n4624) );
  CIVX2 U5558 ( .A(\reg_mem[23][20] ), .Z(n4623) );
  CMXI2X1 U5559 ( .A0(n4626), .A1(n4625), .S(net87624), .Z(n4627) );
  CIVX2 U5560 ( .A(\reg_mem[24][20] ), .Z(n4630) );
  CIVX2 U5561 ( .A(\reg_mem[25][20] ), .Z(n4629) );
  CMXI2X1 U5562 ( .A0(n4630), .A1(n4629), .S(net87797), .Z(n4634) );
  CIVX2 U5563 ( .A(\reg_mem[26][20] ), .Z(n4632) );
  CIVX2 U5564 ( .A(\reg_mem[27][20] ), .Z(n4631) );
  CMXI2X1 U5565 ( .A0(n4632), .A1(n4631), .S(net87800), .Z(n4633) );
  CMXI2X1 U5566 ( .A0(n4634), .A1(n4633), .S(net87631), .Z(n4642) );
  CIVX2 U5567 ( .A(\reg_mem[28][20] ), .Z(n4636) );
  CIVX2 U5568 ( .A(\reg_mem[29][20] ), .Z(n4635) );
  CIVX2 U5569 ( .A(\reg_mem[30][20] ), .Z(n4638) );
  CIVX2 U5570 ( .A(\reg_mem[31][20] ), .Z(n4637) );
  CMXI2X1 U5571 ( .A0(n4638), .A1(n4637), .S(net87793), .Z(n4639) );
  CMXI2X1 U5572 ( .A0(n4640), .A1(n4639), .S(net87628), .Z(n4641) );
  CMXI2X1 U5573 ( .A0(n4642), .A1(n4641), .S(net87730), .Z(n4643) );
  CIVX2 U5574 ( .A(\reg_mem[0][21] ), .Z(n4648) );
  CMXI2X1 U5575 ( .A0(n4648), .A1(n4647), .S(net87799), .Z(n4652) );
  CIVX2 U5576 ( .A(\reg_mem[2][21] ), .Z(n4650) );
  CMXI2X1 U5577 ( .A0(n4650), .A1(n4649), .S(net87798), .Z(n4651) );
  CMXI2X1 U5578 ( .A0(n4652), .A1(n4651), .S(net87635), .Z(n4660) );
  CIVX2 U5579 ( .A(\reg_mem[4][21] ), .Z(n4654) );
  CMXI2X1 U5580 ( .A0(n4654), .A1(n4653), .S(net87802), .Z(n4658) );
  CIVX2 U5581 ( .A(\reg_mem[6][21] ), .Z(n4656) );
  CMXI2X1 U5582 ( .A0(n4656), .A1(n4655), .S(net87807), .Z(n4657) );
  CMXI2X1 U5583 ( .A0(n4658), .A1(n4657), .S(net87634), .Z(n4659) );
  CMXI2X1 U5584 ( .A0(n4660), .A1(n4659), .S(net87710), .Z(n4676) );
  CMXI2X1 U5585 ( .A0(n4662), .A1(n4661), .S(net87802), .Z(n4666) );
  CMXI2X1 U5586 ( .A0(n4664), .A1(n4663), .S(net87794), .Z(n4665) );
  CMXI2X1 U5587 ( .A0(n4666), .A1(n4665), .S(net87626), .Z(n4674) );
  CMXI2X1 U5588 ( .A0(n4668), .A1(n4667), .S(net87794), .Z(n4672) );
  CMXI2X1 U5589 ( .A0(n4670), .A1(n4669), .S(net87802), .Z(n4671) );
  CMXI2X1 U5590 ( .A0(n4672), .A1(n4671), .S(net87639), .Z(n4673) );
  CMXI2X1 U5591 ( .A0(n4674), .A1(n4673), .S(net87718), .Z(n4675) );
  CMXI2X1 U5592 ( .A0(n4676), .A1(n4675), .S(net82865), .Z(n4708) );
  CIVX2 U5593 ( .A(\reg_mem[16][21] ), .Z(n4678) );
  CMXI2X1 U5594 ( .A0(n4678), .A1(n4677), .S(net87793), .Z(n4682) );
  CIVX2 U5595 ( .A(\reg_mem[18][21] ), .Z(n4680) );
  CMXI2X1 U5596 ( .A0(n4680), .A1(n4679), .S(net87794), .Z(n4681) );
  CMXI2X1 U5597 ( .A0(n4682), .A1(n4681), .S(net87636), .Z(n4690) );
  CIVX2 U5598 ( .A(\reg_mem[20][21] ), .Z(n4684) );
  CMXI2X1 U5599 ( .A0(n4684), .A1(n4683), .S(net87802), .Z(n4688) );
  CIVX2 U5600 ( .A(\reg_mem[22][21] ), .Z(n4686) );
  CMXI2X1 U5601 ( .A0(n4686), .A1(n4685), .S(net87799), .Z(n4687) );
  CMXI2X1 U5602 ( .A0(n4690), .A1(n4689), .S(net87727), .Z(n4706) );
  CMXI2X1 U5603 ( .A0(n4692), .A1(n4691), .S(net87807), .Z(n4696) );
  CMXI2X1 U5604 ( .A0(n4694), .A1(n4693), .S(net87806), .Z(n4695) );
  CMXI2X1 U5605 ( .A0(n4696), .A1(n4695), .S(net87623), .Z(n4704) );
  CMXI2X1 U5606 ( .A0(n4698), .A1(n4697), .S(net87793), .Z(n4702) );
  CMXI2X1 U5607 ( .A0(n4700), .A1(n4699), .S(net87806), .Z(n4701) );
  CMXI2X1 U5608 ( .A0(n4702), .A1(n4701), .S(net87636), .Z(n4703) );
  CMXI2X1 U5609 ( .A0(n4704), .A1(n4703), .S(net87706), .Z(n4705) );
  CMXI2X1 U5610 ( .A0(n4706), .A1(n4705), .S(net82865), .Z(n4707) );
  CMXI2X1 U5611 ( .A0(n4708), .A1(n4707), .S(net86657), .Z(N211) );
  CMXI2X1 U5612 ( .A0(n4710), .A1(n4709), .S(net87798), .Z(n4714) );
  CMXI2X1 U5613 ( .A0(n4712), .A1(n4711), .S(net87806), .Z(n4713) );
  CMXI2X1 U5614 ( .A0(n4714), .A1(n4713), .S(net87634), .Z(n4722) );
  CMXI2X1 U5615 ( .A0(n4716), .A1(n4715), .S(net87809), .Z(n4720) );
  CMXI2X1 U5616 ( .A0(n4718), .A1(n4717), .S(net87806), .Z(n4719) );
  CMXI2X1 U5617 ( .A0(n4720), .A1(n4719), .S(net87633), .Z(n4721) );
  CMXI2X1 U5618 ( .A0(n4722), .A1(n4721), .S(net87709), .Z(n4738) );
  CMXI2X1 U5619 ( .A0(n4724), .A1(n4723), .S(net87798), .Z(n4728) );
  CMXI2X1 U5620 ( .A0(n4726), .A1(n4725), .S(net87793), .Z(n4727) );
  CMXI2X1 U5621 ( .A0(n4728), .A1(n4727), .S(net87625), .Z(n4736) );
  CMXI2X1 U5622 ( .A0(n4730), .A1(n4729), .S(net87791), .Z(n4734) );
  CMXI2X1 U5623 ( .A0(n4732), .A1(n4731), .S(net87798), .Z(n4733) );
  CMXI2X1 U5624 ( .A0(n4734), .A1(n4733), .S(net87627), .Z(n4735) );
  CMXI2X1 U5625 ( .A0(n4736), .A1(n4735), .S(net87717), .Z(n4737) );
  CMXI2X1 U5626 ( .A0(n4738), .A1(n4737), .S(net82865), .Z(n4770) );
  CMXI2X1 U5627 ( .A0(n4740), .A1(n4739), .S(net87795), .Z(n4744) );
  CMXI2X1 U5628 ( .A0(n4742), .A1(n4741), .S(net87807), .Z(n4743) );
  CMXI2X1 U5629 ( .A0(n4746), .A1(n4745), .S(net87798), .Z(n4750) );
  CMXI2X1 U5630 ( .A0(n4748), .A1(n4747), .S(net87793), .Z(n4749) );
  CMXI2X1 U5631 ( .A0(n4750), .A1(n4749), .S(net87642), .Z(n4751) );
  CMXI2X1 U5632 ( .A0(n4752), .A1(n4751), .S(net87720), .Z(n4768) );
  CMXI2X1 U5633 ( .A0(n4754), .A1(n4753), .S(net87809), .Z(n4758) );
  CMXI2X1 U5634 ( .A0(n4756), .A1(n4755), .S(net87806), .Z(n4757) );
  CMXI2X1 U5635 ( .A0(n4758), .A1(n4757), .S(net87630), .Z(n4766) );
  CMXI2X1 U5636 ( .A0(n4760), .A1(n4759), .S(net87793), .Z(n4764) );
  CMXI2X1 U5637 ( .A0(n4762), .A1(n4761), .S(net87806), .Z(n4763) );
  CMXI2X1 U5638 ( .A0(n4764), .A1(n4763), .S(net87627), .Z(n4765) );
  CMXI2X1 U5639 ( .A0(n4766), .A1(n4765), .S(net87728), .Z(n4767) );
  CMXI2X1 U5640 ( .A0(n4768), .A1(n4767), .S(net82865), .Z(n4769) );
  CMXI2X1 U5641 ( .A0(n4770), .A1(n4769), .S(net86657), .Z(N210) );
  CMXI2X1 U5642 ( .A0(n4772), .A1(n4771), .S(net87639), .Z(n4778) );
  CIVX2 U5643 ( .A(\reg_mem[6][23] ), .Z(n4774) );
  CIVX2 U5644 ( .A(\reg_mem[7][23] ), .Z(n4773) );
  CMXI2X1 U5645 ( .A0(n4774), .A1(n4773), .S(net87793), .Z(n4775) );
  CMXI2X1 U5646 ( .A0(n4776), .A1(n4775), .S(net87637), .Z(n4777) );
  CMXI2X1 U5647 ( .A0(n4778), .A1(n4777), .S(net87722), .Z(n4788) );
  CMXI2X1 U5648 ( .A0(n4780), .A1(n4779), .S(net87639), .Z(n4786) );
  CIVX2 U5649 ( .A(\reg_mem[14][23] ), .Z(n4782) );
  CIVX2 U5650 ( .A(\reg_mem[15][23] ), .Z(n4781) );
  CMXI2X1 U5651 ( .A0(n4782), .A1(n4781), .S(net87803), .Z(n4783) );
  CMXI2X1 U5652 ( .A0(n4784), .A1(n4783), .S(net87629), .Z(n4785) );
  CMXI2X1 U5653 ( .A0(n4786), .A1(n4785), .S(net87715), .Z(n4787) );
  CMXI2X1 U5654 ( .A0(n4788), .A1(n4787), .S(net82865), .Z(n4814) );
  CMXI2X1 U5655 ( .A0(n4790), .A1(n4789), .S(net87634), .Z(n4796) );
  CIVX2 U5656 ( .A(\reg_mem[22][23] ), .Z(n4792) );
  CMXI2X1 U5657 ( .A0(n4792), .A1(n4791), .S(net87798), .Z(n4793) );
  CMXI2X1 U5658 ( .A0(n4794), .A1(n4793), .S(net87635), .Z(n4795) );
  CMXI2X1 U5659 ( .A0(n4796), .A1(n4795), .S(net87708), .Z(n4812) );
  CIVX2 U5660 ( .A(\reg_mem[24][23] ), .Z(n4798) );
  CIVX2 U5661 ( .A(\reg_mem[25][23] ), .Z(n4797) );
  CMXI2X1 U5662 ( .A0(n4798), .A1(n4797), .S(net87809), .Z(n4802) );
  CIVX2 U5663 ( .A(\reg_mem[26][23] ), .Z(n4800) );
  CIVX2 U5664 ( .A(\reg_mem[27][23] ), .Z(n4799) );
  CMXI2X1 U5665 ( .A0(n4800), .A1(n4799), .S(net87798), .Z(n4801) );
  CMXI2X1 U5666 ( .A0(n4802), .A1(n4801), .S(net87624), .Z(n4810) );
  CIVX2 U5667 ( .A(\reg_mem[28][23] ), .Z(n4804) );
  CIVX2 U5668 ( .A(\reg_mem[29][23] ), .Z(n4803) );
  CMXI2X1 U5669 ( .A0(n4804), .A1(n4803), .S(net87800), .Z(n4808) );
  CIVX2 U5670 ( .A(\reg_mem[30][23] ), .Z(n4806) );
  CIVX2 U5671 ( .A(\reg_mem[31][23] ), .Z(n4805) );
  CMXI2X1 U5672 ( .A0(n4806), .A1(n4805), .S(net87804), .Z(n4807) );
  CMXI2X1 U5673 ( .A0(n4808), .A1(n4807), .S(net87624), .Z(n4809) );
  CMXI2X1 U5674 ( .A0(n4810), .A1(n4809), .S(net87716), .Z(n4811) );
  CMXI2X1 U5675 ( .A0(n4812), .A1(n4811), .S(net82865), .Z(n4813) );
  CIVX2 U5676 ( .A(\reg_mem[6][24] ), .Z(n4818) );
  CIVX2 U5677 ( .A(\reg_mem[7][24] ), .Z(n4817) );
  CMXI2X1 U5678 ( .A0(n4818), .A1(n4817), .S(net87797), .Z(n4819) );
  CMXI2X1 U5679 ( .A0(n4820), .A1(n4819), .S(net87635), .Z(n4821) );
  CMXI2X1 U5680 ( .A0(n4822), .A1(n4821), .S(net87714), .Z(n4832) );
  CIVX2 U5681 ( .A(\reg_mem[14][24] ), .Z(n4826) );
  CIVX2 U5682 ( .A(\reg_mem[15][24] ), .Z(n4825) );
  CMXI2X1 U5683 ( .A0(n4826), .A1(n4825), .S(net87794), .Z(n4827) );
  CMXI2X1 U5684 ( .A0(n4830), .A1(n4829), .S(net87714), .Z(n4831) );
  CMXI2X1 U5685 ( .A0(n4832), .A1(n4831), .S(net82867), .Z(n4858) );
  CIVX2 U5686 ( .A(\reg_mem[22][24] ), .Z(n4836) );
  CIVX2 U5687 ( .A(\reg_mem[23][24] ), .Z(n4835) );
  CMXI2X1 U5688 ( .A0(n4838), .A1(n4837), .S(net87632), .Z(n4839) );
  CMXI2X1 U5689 ( .A0(n4840), .A1(n4839), .S(net87724), .Z(n4856) );
  CIVX2 U5690 ( .A(\reg_mem[24][24] ), .Z(n4842) );
  CIVX2 U5691 ( .A(\reg_mem[25][24] ), .Z(n4841) );
  CMXI2X1 U5692 ( .A0(n4842), .A1(n4841), .S(net87798), .Z(n4846) );
  CIVX2 U5693 ( .A(\reg_mem[26][24] ), .Z(n4844) );
  CIVX2 U5694 ( .A(\reg_mem[27][24] ), .Z(n4843) );
  CMXI2X1 U5695 ( .A0(n4844), .A1(n4843), .S(net87809), .Z(n4845) );
  CIVX2 U5696 ( .A(\reg_mem[28][24] ), .Z(n4848) );
  CIVX2 U5697 ( .A(\reg_mem[29][24] ), .Z(n4847) );
  CMXI2X1 U5698 ( .A0(n4848), .A1(n4847), .S(net87800), .Z(n4852) );
  CIVX2 U5699 ( .A(\reg_mem[30][24] ), .Z(n4850) );
  CIVX2 U5700 ( .A(\reg_mem[31][24] ), .Z(n4849) );
  CMXI2X1 U5701 ( .A0(n4850), .A1(n4849), .S(net87806), .Z(n4851) );
  CMXI2X1 U5702 ( .A0(n4854), .A1(n4853), .S(net87715), .Z(n4855) );
  CMXI2X1 U5703 ( .A0(n4860), .A1(n4859), .S(net87793), .Z(n4864) );
  CMXI2X1 U5704 ( .A0(n4862), .A1(n4861), .S(net87797), .Z(n4863) );
  CMXI2X1 U5705 ( .A0(n4864), .A1(n4863), .S(net87633), .Z(n4872) );
  CMXI2X1 U5706 ( .A0(n4866), .A1(n4865), .S(net87797), .Z(n4870) );
  CMXI2X1 U5707 ( .A0(n4870), .A1(n4869), .S(net87632), .Z(n4871) );
  CMXI2X1 U5708 ( .A0(n4872), .A1(n4871), .S(net87708), .Z(n4888) );
  CMXI2X1 U5709 ( .A0(n4874), .A1(n4873), .S(net87800), .Z(n4878) );
  CMXI2X1 U5710 ( .A0(n4876), .A1(n4875), .S(net87793), .Z(n4877) );
  CMXI2X1 U5711 ( .A0(n4878), .A1(n4877), .S(net87624), .Z(n4886) );
  CMXI2X1 U5712 ( .A0(n4882), .A1(n4881), .S(net87807), .Z(n4883) );
  CMXI2X1 U5713 ( .A0(n4884), .A1(n4883), .S(net87626), .Z(n4885) );
  CMXI2X1 U5714 ( .A0(n4886), .A1(n4885), .S(net87716), .Z(n4887) );
  CMXI2X1 U5715 ( .A0(n4888), .A1(n4887), .S(net82867), .Z(n4920) );
  CMXI2X1 U5716 ( .A0(n4890), .A1(n4889), .S(net87800), .Z(n4894) );
  CMXI2X1 U5717 ( .A0(n4892), .A1(n4891), .S(net87804), .Z(n4893) );
  CMXI2X1 U5718 ( .A0(n4894), .A1(n4893), .S(net87640), .Z(n4902) );
  CMXI2X1 U5719 ( .A0(n4896), .A1(n4895), .S(net87803), .Z(n4900) );
  CMXI2X1 U5720 ( .A0(n4898), .A1(n4897), .S(net87803), .Z(n4899) );
  CMXI2X1 U5721 ( .A0(n4900), .A1(n4899), .S(net87642), .Z(n4901) );
  CMXI2X1 U5722 ( .A0(n4902), .A1(n4901), .S(net87706), .Z(n4918) );
  CMXI2X1 U5723 ( .A0(n4904), .A1(n4903), .S(net87802), .Z(n4908) );
  CMXI2X1 U5724 ( .A0(n4906), .A1(n4905), .S(net87794), .Z(n4907) );
  CMXI2X1 U5725 ( .A0(n4908), .A1(n4907), .S(net87629), .Z(n4916) );
  CMXI2X1 U5726 ( .A0(n4910), .A1(n4909), .S(net87791), .Z(n4914) );
  CMXI2X1 U5727 ( .A0(n4912), .A1(n4911), .S(net87800), .Z(n4913) );
  CMXI2X1 U5728 ( .A0(n4914), .A1(n4913), .S(net87623), .Z(n4915) );
  CMXI2X1 U5729 ( .A0(n4916), .A1(n4915), .S(net87727), .Z(n4917) );
  CMXI2X1 U5730 ( .A0(n4918), .A1(n4917), .S(net82867), .Z(n4919) );
  CMXI2X1 U5731 ( .A0(n4920), .A1(n4919), .S(net86657), .Z(N207) );
  CMXI2X1 U5732 ( .A0(n4922), .A1(n4921), .S(net87797), .Z(n4926) );
  CMXI2X1 U5733 ( .A0(n4924), .A1(n4923), .S(net87794), .Z(n4925) );
  CMXI2X1 U5734 ( .A0(n4926), .A1(n4925), .S(net87631), .Z(n4934) );
  CMXI2X1 U5735 ( .A0(n4928), .A1(n4927), .S(net87795), .Z(n4932) );
  CMXI2X1 U5736 ( .A0(n4930), .A1(n4929), .S(net87809), .Z(n4931) );
  CMXI2X1 U5737 ( .A0(n4932), .A1(n4931), .S(net87638), .Z(n4933) );
  CMXI2X1 U5738 ( .A0(n4934), .A1(n4933), .S(net87718), .Z(n4950) );
  CMXI2X1 U5739 ( .A0(n4936), .A1(n4935), .S(net87806), .Z(n4940) );
  CMXI2X1 U5740 ( .A0(n4938), .A1(n4937), .S(net87804), .Z(n4939) );
  CMXI2X1 U5741 ( .A0(n4940), .A1(n4939), .S(net87630), .Z(n4948) );
  CMXI2X1 U5742 ( .A0(n4942), .A1(n4941), .S(net87793), .Z(n4946) );
  CMXI2X1 U5743 ( .A0(n4944), .A1(n4943), .S(net87804), .Z(n4945) );
  CMXI2X1 U5744 ( .A0(n4946), .A1(n4945), .S(net87623), .Z(n4947) );
  CMXI2X1 U5745 ( .A0(n4948), .A1(n4947), .S(net87715), .Z(n4949) );
  CMXI2X1 U5746 ( .A0(n4950), .A1(n4949), .S(net82867), .Z(n4982) );
  CMXI2X1 U5747 ( .A0(n4952), .A1(n4951), .S(net87791), .Z(n4956) );
  CMXI2X1 U5748 ( .A0(n4954), .A1(n4953), .S(net87803), .Z(n4955) );
  CMXI2X1 U5749 ( .A0(n4956), .A1(n4955), .S(net87639), .Z(n4964) );
  CMXI2X1 U5750 ( .A0(n4958), .A1(n4957), .S(net87803), .Z(n4962) );
  CMXI2X1 U5751 ( .A0(n4960), .A1(n4959), .S(net87803), .Z(n4961) );
  CMXI2X1 U5752 ( .A0(n4964), .A1(n4963), .S(net87705), .Z(n4980) );
  CMXI2X1 U5753 ( .A0(n4966), .A1(n4965), .S(net87809), .Z(n4970) );
  CMXI2X1 U5754 ( .A0(n4968), .A1(n4967), .S(net87803), .Z(n4969) );
  CMXI2X1 U5755 ( .A0(n4970), .A1(n4969), .S(net87628), .Z(n4978) );
  CMXI2X1 U5756 ( .A0(n4972), .A1(n4971), .S(net87797), .Z(n4976) );
  CMXI2X1 U5757 ( .A0(n4974), .A1(n4973), .S(net87809), .Z(n4975) );
  CMXI2X1 U5758 ( .A0(n4976), .A1(n4975), .S(net87639), .Z(n4977) );
  CMXI2X1 U5759 ( .A0(n4978), .A1(n4977), .S(net87725), .Z(n4979) );
  CMXI2X1 U5760 ( .A0(n4980), .A1(n4979), .S(net82867), .Z(n4981) );
  CMXI2X1 U5761 ( .A0(n4982), .A1(n4981), .S(net86657), .Z(N206) );
  CMXI2X1 U5762 ( .A0(n4986), .A1(n4985), .S(net87706), .Z(n4996) );
  CIVX2 U5763 ( .A(\reg_mem[14][27] ), .Z(n4990) );
  CIVX2 U5764 ( .A(\reg_mem[15][27] ), .Z(n4989) );
  CMXI2X1 U5765 ( .A0(n4990), .A1(n4989), .S(net87807), .Z(n4991) );
  CMXI2X1 U5766 ( .A0(n4998), .A1(n4997), .S(net87635), .Z(n5004) );
  CIVX2 U5767 ( .A(\reg_mem[22][27] ), .Z(n5000) );
  CIVX2 U5768 ( .A(\reg_mem[23][27] ), .Z(n4999) );
  CMXI2X1 U5769 ( .A0(n5000), .A1(n4999), .S(net87804), .Z(n5001) );
  CMXI2X1 U5770 ( .A0(n5004), .A1(n5003), .S(net87704), .Z(n5020) );
  CIVX2 U5771 ( .A(\reg_mem[24][27] ), .Z(n5006) );
  CIVX2 U5772 ( .A(\reg_mem[25][27] ), .Z(n5005) );
  CMXI2X1 U5773 ( .A0(n5006), .A1(n5005), .S(net87798), .Z(n5010) );
  CIVX2 U5774 ( .A(\reg_mem[26][27] ), .Z(n5008) );
  CIVX2 U5775 ( .A(\reg_mem[27][27] ), .Z(n5007) );
  CMXI2X1 U5776 ( .A0(n5008), .A1(n5007), .S(net87807), .Z(n5009) );
  CMXI2X1 U5777 ( .A0(n5010), .A1(n5009), .S(net87625), .Z(n5018) );
  CIVX2 U5778 ( .A(\reg_mem[28][27] ), .Z(n5012) );
  CIVX2 U5779 ( .A(\reg_mem[29][27] ), .Z(n5011) );
  CMXI2X1 U5780 ( .A0(n5012), .A1(n5011), .S(net87791), .Z(n5016) );
  CIVX2 U5781 ( .A(\reg_mem[30][27] ), .Z(n5014) );
  CIVX2 U5782 ( .A(\reg_mem[31][27] ), .Z(n5013) );
  CMXI2X1 U5783 ( .A0(n5014), .A1(n5013), .S(net87793), .Z(n5015) );
  CMXI2X1 U5784 ( .A0(n5016), .A1(n5015), .S(net87635), .Z(n5017) );
  CMXI2X1 U5785 ( .A0(n5018), .A1(n5017), .S(net87725), .Z(n5019) );
  CIVX2 U5786 ( .A(\reg_mem[6][28] ), .Z(n5024) );
  CIVX2 U5787 ( .A(\reg_mem[7][28] ), .Z(n5023) );
  CMXI2X1 U5788 ( .A0(n5024), .A1(n5023), .S(net87809), .Z(n5025) );
  CMXI2X1 U5789 ( .A0(n5026), .A1(n5025), .S(net87632), .Z(n5027) );
  CMXI2X1 U5790 ( .A0(n5028), .A1(n5027), .S(net87710), .Z(n5038) );
  CMXI2X1 U5791 ( .A0(n5030), .A1(n5029), .S(net87636), .Z(n5036) );
  CIVX2 U5792 ( .A(\reg_mem[14][28] ), .Z(n5032) );
  CIVX2 U5793 ( .A(\reg_mem[15][28] ), .Z(n5031) );
  CMXI2X1 U5794 ( .A0(n5032), .A1(n5031), .S(net87802), .Z(n5033) );
  CMXI2X1 U5795 ( .A0(n5034), .A1(n5033), .S(net87628), .Z(n5035) );
  CMXI2X1 U5796 ( .A0(n5036), .A1(n5035), .S(net87709), .Z(n5037) );
  CMXI2X1 U5797 ( .A0(n5038), .A1(n5037), .S(net82867), .Z(n5064) );
  CMXI2X1 U5798 ( .A0(n5040), .A1(n5039), .S(net87633), .Z(n5046) );
  CIVX2 U5799 ( .A(\reg_mem[22][28] ), .Z(n5042) );
  CIVX2 U5800 ( .A(\reg_mem[23][28] ), .Z(n5041) );
  CMXI2X1 U5801 ( .A0(n5042), .A1(n5041), .S(net87809), .Z(n5043) );
  CMXI2X1 U5802 ( .A0(n5044), .A1(n5043), .S(net87634), .Z(n5045) );
  CMXI2X1 U5803 ( .A0(n5046), .A1(n5045), .S(net87720), .Z(n5062) );
  CIVX2 U5804 ( .A(\reg_mem[24][28] ), .Z(n5048) );
  CIVX2 U5805 ( .A(\reg_mem[25][28] ), .Z(n5047) );
  CMXI2X1 U5806 ( .A0(n5048), .A1(n5047), .S(net87799), .Z(n5052) );
  CIVX2 U5807 ( .A(\reg_mem[26][28] ), .Z(n5050) );
  CIVX2 U5808 ( .A(\reg_mem[27][28] ), .Z(n5049) );
  CMXI2X1 U5809 ( .A0(n5050), .A1(n5049), .S(net87798), .Z(n5051) );
  CMXI2X1 U5810 ( .A0(n5052), .A1(n5051), .S(net87623), .Z(n5060) );
  CIVX2 U5811 ( .A(\reg_mem[28][28] ), .Z(n5054) );
  CIVX2 U5812 ( .A(\reg_mem[29][28] ), .Z(n5053) );
  CMXI2X1 U5813 ( .A0(n5054), .A1(n5053), .S(net87791), .Z(n5058) );
  CIVX2 U5814 ( .A(\reg_mem[30][28] ), .Z(n5056) );
  CIVX2 U5815 ( .A(\reg_mem[31][28] ), .Z(n5055) );
  CMXI2X1 U5816 ( .A0(n5056), .A1(n5055), .S(net87809), .Z(n5057) );
  CMXI2X1 U5817 ( .A0(n5058), .A1(n5057), .S(net87623), .Z(n5059) );
  CMXI2X1 U5818 ( .A0(n5060), .A1(n5059), .S(net87714), .Z(n5061) );
  CMXI2X1 U5819 ( .A0(n5062), .A1(n5061), .S(net82867), .Z(n5063) );
  CIVX2 U5820 ( .A(\reg_mem[2][29] ), .Z(n5066) );
  CIVX2 U5821 ( .A(\reg_mem[3][29] ), .Z(n5065) );
  CMXI2X1 U5822 ( .A0(n5066), .A1(n5065), .S(net87802), .Z(n5067) );
  CMXI2X1 U5823 ( .A0(n5068), .A1(n5067), .S(net87638), .Z(n5076) );
  CIVX2 U5824 ( .A(\reg_mem[4][29] ), .Z(n5070) );
  CIVX2 U5825 ( .A(\reg_mem[5][29] ), .Z(n5069) );
  CMXI2X1 U5826 ( .A0(n5070), .A1(n5069), .S(net87806), .Z(n5074) );
  CIVX2 U5827 ( .A(\reg_mem[6][29] ), .Z(n5072) );
  CIVX2 U5828 ( .A(\reg_mem[7][29] ), .Z(n5071) );
  CMXI2X1 U5829 ( .A0(n5072), .A1(n5071), .S(net87800), .Z(n5073) );
  CMXI2X1 U5830 ( .A0(n5074), .A1(n5073), .S(net87636), .Z(n5075) );
  CMXI2X1 U5831 ( .A0(n5076), .A1(n5075), .S(net87710), .Z(n5084) );
  CIVX2 U5832 ( .A(\reg_mem[14][29] ), .Z(n5078) );
  CIVX2 U5833 ( .A(\reg_mem[15][29] ), .Z(n5077) );
  CMXI2X1 U5834 ( .A0(n5078), .A1(n5077), .S(net87802), .Z(n5079) );
  CMXI2X1 U5835 ( .A0(n5080), .A1(n5079), .S(net87630), .Z(n5081) );
  CMXI2X1 U5836 ( .A0(n5082), .A1(n5081), .S(net87728), .Z(n5083) );
  CMXI2X1 U5837 ( .A0(n5084), .A1(n5083), .S(net82867), .Z(n5114) );
  CIVX2 U5838 ( .A(\reg_mem[18][29] ), .Z(n5086) );
  CIVX2 U5839 ( .A(\reg_mem[19][29] ), .Z(n5085) );
  CMXI2X1 U5840 ( .A0(n5086), .A1(n5085), .S(net87797), .Z(n5087) );
  CMXI2X1 U5841 ( .A0(n5088), .A1(n5087), .S(net87632), .Z(n5096) );
  CIVX2 U5842 ( .A(\reg_mem[20][29] ), .Z(n5090) );
  CIVX2 U5843 ( .A(\reg_mem[21][29] ), .Z(n5089) );
  CMXI2X1 U5844 ( .A0(n5090), .A1(n5089), .S(net87803), .Z(n5094) );
  CIVX2 U5845 ( .A(\reg_mem[22][29] ), .Z(n5092) );
  CIVX2 U5846 ( .A(\reg_mem[23][29] ), .Z(n5091) );
  CMXI2X1 U5847 ( .A0(n5092), .A1(n5091), .S(net87806), .Z(n5093) );
  CMXI2X1 U5848 ( .A0(n5094), .A1(n5093), .S(net87633), .Z(n5095) );
  CMXI2X1 U5849 ( .A0(n5096), .A1(n5095), .S(net87719), .Z(n5112) );
  CIVX2 U5850 ( .A(\reg_mem[24][29] ), .Z(n5098) );
  CIVX2 U5851 ( .A(\reg_mem[25][29] ), .Z(n5097) );
  CMXI2X1 U5852 ( .A0(n5098), .A1(n5097), .S(net87798), .Z(n5102) );
  CIVX2 U5853 ( .A(\reg_mem[26][29] ), .Z(n5100) );
  CIVX2 U5854 ( .A(\reg_mem[27][29] ), .Z(n5099) );
  CMXI2X1 U5855 ( .A0(n5100), .A1(n5099), .S(net87800), .Z(n5101) );
  CMXI2X1 U5856 ( .A0(n5102), .A1(n5101), .S(net87642), .Z(n5110) );
  CIVX2 U5857 ( .A(\reg_mem[28][29] ), .Z(n5104) );
  CIVX2 U5858 ( .A(\reg_mem[29][29] ), .Z(n5103) );
  CIVX2 U5859 ( .A(\reg_mem[30][29] ), .Z(n5106) );
  CIVX2 U5860 ( .A(\reg_mem[31][29] ), .Z(n5105) );
  CMXI2X1 U5861 ( .A0(n5106), .A1(n5105), .S(net87791), .Z(n5107) );
  CMXI2X1 U5862 ( .A0(n5108), .A1(n5107), .S(net87642), .Z(n5109) );
  CMXI2X1 U5863 ( .A0(n5110), .A1(n5109), .S(net87730), .Z(n5111) );
  CMXI2X1 U5864 ( .A0(n5112), .A1(n5111), .S(net82867), .Z(n5113) );
  CMXI2X1 U5865 ( .A0(n5114), .A1(n5113), .S(net86657), .Z(N203) );
  CMXI2X1 U5866 ( .A0(n5116), .A1(n5115), .S(net87635), .Z(n5122) );
  CIVX2 U5867 ( .A(\reg_mem[6][30] ), .Z(n5118) );
  CIVX2 U5868 ( .A(\reg_mem[7][30] ), .Z(n5117) );
  CMXI2X1 U5869 ( .A0(n5118), .A1(n5117), .S(net87794), .Z(n5119) );
  CMXI2X1 U5870 ( .A0(n5120), .A1(n5119), .S(net87627), .Z(n5121) );
  CMXI2X1 U5871 ( .A0(n5122), .A1(n5121), .S(net87719), .Z(n5132) );
  CMXI2X1 U5872 ( .A0(n5124), .A1(n5123), .S(net87630), .Z(n5130) );
  CIVX2 U5873 ( .A(\reg_mem[14][30] ), .Z(n5126) );
  CIVX2 U5874 ( .A(\reg_mem[15][30] ), .Z(n5125) );
  CMXI2X1 U5875 ( .A0(n5126), .A1(n5125), .S(net87803), .Z(n5127) );
  CMXI2X1 U5876 ( .A0(n5128), .A1(n5127), .S(net87631), .Z(n5129) );
  CMXI2X1 U5877 ( .A0(n5130), .A1(n5129), .S(net87709), .Z(n5131) );
  CMXI2X1 U5878 ( .A0(n5134), .A1(n5133), .S(net87630), .Z(n5140) );
  CIVX2 U5879 ( .A(\reg_mem[22][30] ), .Z(n5136) );
  CIVX2 U5880 ( .A(\reg_mem[23][30] ), .Z(n5135) );
  CMXI2X1 U5881 ( .A0(n5136), .A1(n5135), .S(net87809), .Z(n5137) );
  CMXI2X1 U5882 ( .A0(n5138), .A1(n5137), .S(net87637), .Z(n5139) );
  CMXI2X1 U5883 ( .A0(n5140), .A1(n5139), .S(net87718), .Z(n5156) );
  CIVX2 U5884 ( .A(\reg_mem[24][30] ), .Z(n5142) );
  CIVX2 U5885 ( .A(\reg_mem[25][30] ), .Z(n5141) );
  CMXI2X1 U5886 ( .A0(n5142), .A1(n5141), .S(net87804), .Z(n5146) );
  CIVX2 U5887 ( .A(\reg_mem[26][30] ), .Z(n5144) );
  CIVX2 U5888 ( .A(\reg_mem[27][30] ), .Z(n5143) );
  CMXI2X1 U5889 ( .A0(n5144), .A1(n5143), .S(net87791), .Z(n5145) );
  CMXI2X1 U5890 ( .A0(n5146), .A1(n5145), .S(net87640), .Z(n5154) );
  CIVX2 U5891 ( .A(\reg_mem[28][30] ), .Z(n5148) );
  CIVX2 U5892 ( .A(\reg_mem[29][30] ), .Z(n5147) );
  CMXI2X1 U5893 ( .A0(n5148), .A1(n5147), .S(net87806), .Z(n5152) );
  CIVX2 U5894 ( .A(\reg_mem[30][30] ), .Z(n5150) );
  CIVX2 U5895 ( .A(\reg_mem[31][30] ), .Z(n5149) );
  CMXI2X1 U5896 ( .A0(n5150), .A1(n5149), .S(net87806), .Z(n5151) );
  CMXI2X1 U5897 ( .A0(n5152), .A1(n5151), .S(net87640), .Z(n5153) );
  CMXI2X1 U5898 ( .A0(n5154), .A1(n5153), .S(net87719), .Z(n5155) );
  CMXI2X1 U5899 ( .A0(n5156), .A1(n5155), .S(net82869), .Z(n5157) );
  CIVX2 U5900 ( .A(\reg_mem[1][31] ), .Z(n5159) );
  CMXI2X1 U5901 ( .A0(n5160), .A1(n5159), .S(net87799), .Z(n5164) );
  CIVX2 U5902 ( .A(\reg_mem[3][31] ), .Z(n5161) );
  CMXI2X1 U5903 ( .A0(n5162), .A1(n5161), .S(net87799), .Z(n5163) );
  CMXI2X1 U5904 ( .A0(n5164), .A1(n5163), .S(net87629), .Z(n5172) );
  CIVX2 U5905 ( .A(\reg_mem[5][31] ), .Z(n5165) );
  CMXI2X1 U5906 ( .A0(n5166), .A1(n5165), .S(net87803), .Z(n5170) );
  CIVX2 U5907 ( .A(\reg_mem[7][31] ), .Z(n5167) );
  CMXI2X1 U5908 ( .A0(n5168), .A1(n5167), .S(net87795), .Z(n5169) );
  CMXI2X1 U5909 ( .A0(n5170), .A1(n5169), .S(net87630), .Z(n5171) );
  CMXI2X1 U5910 ( .A0(n5172), .A1(n5171), .S(net87708), .Z(n5182) );
  CIVX2 U5911 ( .A(\reg_mem[14][31] ), .Z(n5176) );
  CIVX2 U5912 ( .A(\reg_mem[15][31] ), .Z(n5175) );
  CMXI2X1 U5913 ( .A0(n5176), .A1(n5175), .S(net87793), .Z(n5177) );
  CMXI2X1 U5914 ( .A0(n5178), .A1(n5177), .S(net87626), .Z(n5179) );
  CMXI2X1 U5915 ( .A0(n5180), .A1(n5179), .S(net87710), .Z(n5181) );
  CMXI2X1 U5916 ( .A0(n5182), .A1(n5181), .S(net82869), .Z(n5214) );
  CIVX2 U5917 ( .A(\reg_mem[17][31] ), .Z(n5183) );
  CMXI2X1 U5918 ( .A0(n5184), .A1(n5183), .S(net87806), .Z(n5188) );
  CIVX2 U5919 ( .A(\reg_mem[19][31] ), .Z(n5185) );
  CMXI2X1 U5920 ( .A0(n5186), .A1(n5185), .S(net87809), .Z(n5187) );
  CMXI2X1 U5921 ( .A0(n5188), .A1(n5187), .S(net87626), .Z(n5196) );
  CIVX2 U5922 ( .A(\reg_mem[21][31] ), .Z(n5189) );
  CMXI2X1 U5923 ( .A0(n5190), .A1(n5189), .S(net87807), .Z(n5194) );
  CIVX2 U5924 ( .A(\reg_mem[23][31] ), .Z(n5191) );
  CMXI2X1 U5925 ( .A0(n5194), .A1(n5193), .S(net87635), .Z(n5195) );
  CMXI2X1 U5926 ( .A0(n5196), .A1(n5195), .S(net87717), .Z(n5212) );
  CIVX2 U5927 ( .A(\reg_mem[24][31] ), .Z(n5198) );
  CIVX2 U5928 ( .A(\reg_mem[25][31] ), .Z(n5197) );
  CMXI2X1 U5929 ( .A0(n5198), .A1(n5197), .S(net87809), .Z(n5202) );
  CIVX2 U5930 ( .A(\reg_mem[26][31] ), .Z(n5200) );
  CIVX2 U5931 ( .A(\reg_mem[27][31] ), .Z(n5199) );
  CMXI2X1 U5932 ( .A0(n5200), .A1(n5199), .S(net87791), .Z(n5201) );
  CIVX2 U5933 ( .A(\reg_mem[28][31] ), .Z(n5204) );
  CIVX2 U5934 ( .A(\reg_mem[29][31] ), .Z(n5203) );
  CMXI2X1 U5935 ( .A0(n5204), .A1(n5203), .S(net87791), .Z(n5208) );
  CIVX2 U5936 ( .A(\reg_mem[30][31] ), .Z(n5206) );
  CIVX2 U5937 ( .A(\reg_mem[31][31] ), .Z(n5205) );
  CMXI2X1 U5938 ( .A0(n5206), .A1(n5205), .S(net87794), .Z(n5207) );
  CMXI2X1 U5939 ( .A0(n5208), .A1(n5207), .S(net87636), .Z(n5209) );
  CMXI2X1 U5940 ( .A0(n5210), .A1(n5209), .S(net87718), .Z(n5211) );
  CMXI2X1 U5941 ( .A0(n5212), .A1(n5211), .S(net82869), .Z(n5213) );
  CIVX2 U5942 ( .A(opcode_ex[0]), .Z(n5241) );
  CND2IX1 U5943 ( .B(net76777), .A(n5235), .Z(immi_val_c[16]) );
  CND2IX1 U5944 ( .B(net76776), .A(n5235), .Z(immi_val_c[17]) );
  CND2IX1 U5945 ( .B(n5228), .A(n5235), .Z(immi_val_c[18]) );
  CND2IX1 U5946 ( .B(n5229), .A(n5235), .Z(immi_val_c[19]) );
  CND2IX1 U5947 ( .B(n5230), .A(n5235), .Z(immi_val_c[20]) );
  CND2IX1 U5948 ( .B(n5231), .A(n5235), .Z(immi_val_c[21]) );
  CND2IX1 U5949 ( .B(n5232), .A(n5235), .Z(immi_val_c[22]) );
  CND2IX1 U5950 ( .B(n5233), .A(n5235), .Z(immi_val_c[23]) );
  CND2IX1 U5951 ( .B(n5234), .A(n5235), .Z(immi_val_c[24]) );
  CND2IX1 U5952 ( .B(n5236), .A(n5235), .Z(immi_val_c[25]) );
  CIVX2 U5953 ( .A(inst_fetch[21]), .Z(n5247) );
  CIVX2 U5954 ( .A(inst_fetch[20]), .Z(n5248) );
  CIVX2 U5955 ( .A(inst_fetch[19]), .Z(n5249) );
  CIVX2 U5956 ( .A(inst_fetch[18]), .Z(n5250) );
  CIVX2 U5957 ( .A(inst_fetch[17]), .Z(n5251) );
  CIVX2 U5958 ( .A(inst_fetch[16]), .Z(n5252) );
  CIVX2 U5959 ( .A(inst_fetch[15]), .Z(n5253) );
  CIVX2 U5960 ( .A(inst_fetch[14]), .Z(n5254) );
  CIVX2 U5961 ( .A(inst_fetch[13]), .Z(n5255) );
  CIVX2 U5962 ( .A(inst_fetch[12]), .Z(n5256) );
  CIVX2 U5963 ( .A(inst_fetch[11]), .Z(n5257) );
  CIVX2 U5964 ( .A(inst_fetch[10]), .Z(n5258) );
  CIVX2 U5965 ( .A(inst_fetch[9]), .Z(n5259) );
  CIVX2 U5966 ( .A(inst_fetch[8]), .Z(n5260) );
  CIVX2 U5967 ( .A(inst_fetch[7]), .Z(n5261) );
  CIVX2 U5968 ( .A(inst_fetch[6]), .Z(n5262) );
  CIVX2 U5969 ( .A(opcode_ex[1]), .Z(n5264) );
  CIVX2 U5970 ( .A(n208), .Z(n5265) );
  CIVX2 U5971 ( .A(n231), .Z(n5266) );
  CIVX2 U5972 ( .A(n229), .Z(n5267) );
  CIVX2 U5973 ( .A(opcode_mem[2]), .Z(n5268) );
endmodule

